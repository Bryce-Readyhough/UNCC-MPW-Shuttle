magic
tech sky130A
<<<<<<< HEAD
timestamp 1606420262
=======
timestamp 1606416959
<< checkpaint >>
rect -4848 -4313 296810 356281
>>>>>>> upstream/master
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4411 -480 4467 240
rect 5009 -480 5065 240
rect 5607 -480 5663 240
rect 6205 -480 6261 240
rect 6803 -480 6859 240
rect 7401 -480 7457 240
rect 7999 -480 8055 240
rect 8597 -480 8653 240
rect 9149 -480 9205 240
rect 9747 -480 9803 240
rect 10345 -480 10401 240
rect 10943 -480 10999 240
rect 11541 -480 11597 240
rect 12139 -480 12195 240
rect 12737 -480 12793 240
rect 13335 -480 13391 240
rect 13933 -480 13989 240
rect 14531 -480 14587 240
rect 15129 -480 15185 240
rect 15727 -480 15783 240
rect 16325 -480 16381 240
rect 16923 -480 16979 240
rect 17475 -480 17531 240
rect 18073 -480 18129 240
rect 18671 -480 18727 240
rect 19269 -480 19325 240
rect 19867 -480 19923 240
rect 20465 -480 20521 240
rect 21063 -480 21119 240
rect 21661 -480 21717 240
rect 22259 -480 22315 240
rect 22857 -480 22913 240
rect 23455 -480 23511 240
rect 24053 -480 24109 240
rect 24651 -480 24707 240
rect 25249 -480 25305 240
rect 25801 -480 25857 240
rect 26399 -480 26455 240
rect 26997 -480 27053 240
rect 27595 -480 27651 240
rect 28193 -480 28249 240
rect 28791 -480 28847 240
rect 29389 -480 29445 240
rect 29987 -480 30043 240
rect 30585 -480 30641 240
rect 31183 -480 31239 240
rect 31781 -480 31837 240
rect 32379 -480 32435 240
rect 32977 -480 33033 240
rect 33575 -480 33631 240
rect 34127 -480 34183 240
rect 34725 -480 34781 240
rect 35323 -480 35379 240
rect 35921 -480 35977 240
rect 36519 -480 36575 240
rect 37117 -480 37173 240
rect 37715 -480 37771 240
rect 38313 -480 38369 240
rect 38911 -480 38967 240
rect 39509 -480 39565 240
rect 40107 -480 40163 240
rect 40705 -480 40761 240
rect 41303 -480 41359 240
rect 41901 -480 41957 240
rect 42453 -480 42509 240
rect 43051 -480 43107 240
rect 43649 -480 43705 240
rect 44247 -480 44303 240
rect 44845 -480 44901 240
rect 45443 -480 45499 240
rect 46041 -480 46097 240
rect 46639 -480 46695 240
rect 47237 -480 47293 240
rect 47835 -480 47891 240
rect 48433 -480 48489 240
rect 49031 -480 49087 240
rect 49629 -480 49685 240
rect 50227 -480 50283 240
rect 50779 -480 50835 240
rect 51377 -480 51433 240
rect 51975 -480 52031 240
rect 52573 -480 52629 240
rect 53171 -480 53227 240
rect 53769 -480 53825 240
rect 54367 -480 54423 240
rect 54965 -480 55021 240
rect 55563 -480 55619 240
rect 56161 -480 56217 240
rect 56759 -480 56815 240
rect 57357 -480 57413 240
rect 57955 -480 58011 240
rect 58553 -480 58609 240
rect 59105 -480 59161 240
rect 59703 -480 59759 240
rect 60301 -480 60357 240
rect 60899 -480 60955 240
rect 61497 -480 61553 240
rect 62095 -480 62151 240
rect 62693 -480 62749 240
rect 63291 -480 63347 240
rect 63889 -480 63945 240
rect 64487 -480 64543 240
rect 65085 -480 65141 240
rect 65683 -480 65739 240
rect 66281 -480 66337 240
rect 66879 -480 66935 240
rect 67431 -480 67487 240
rect 68029 -480 68085 240
rect 68627 -480 68683 240
rect 69225 -480 69281 240
rect 69823 -480 69879 240
rect 70421 -480 70477 240
rect 71019 -480 71075 240
rect 71617 -480 71673 240
rect 72215 -480 72271 240
rect 72813 -480 72869 240
rect 73411 -480 73467 240
rect 74009 -480 74065 240
rect 74607 -480 74663 240
rect 75205 -480 75261 240
rect 75757 -480 75813 240
rect 76355 -480 76411 240
rect 76953 -480 77009 240
rect 77551 -480 77607 240
rect 78149 -480 78205 240
rect 78747 -480 78803 240
rect 79345 -480 79401 240
rect 79943 -480 79999 240
rect 80541 -480 80597 240
rect 81139 -480 81195 240
rect 81737 -480 81793 240
rect 82335 -480 82391 240
rect 82933 -480 82989 240
rect 83531 -480 83587 240
rect 84083 -480 84139 240
rect 84681 -480 84737 240
rect 85279 -480 85335 240
rect 85877 -480 85933 240
rect 86475 -480 86531 240
rect 87073 -480 87129 240
rect 87671 -480 87727 240
rect 88269 -480 88325 240
rect 88867 -480 88923 240
rect 89465 -480 89521 240
rect 90063 -480 90119 240
rect 90661 -480 90717 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92409 -480 92465 240
rect 93007 -480 93063 240
rect 93605 -480 93661 240
rect 94203 -480 94259 240
rect 94801 -480 94857 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98987 -480 99043 240
rect 99585 -480 99641 240
rect 100183 -480 100239 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103127 -480 103183 240
rect 103725 -480 103781 240
rect 104323 -480 104379 240
rect 104921 -480 104977 240
rect 105519 -480 105575 240
rect 106117 -480 106173 240
rect 106715 -480 106771 240
rect 107313 -480 107369 240
rect 107911 -480 107967 240
rect 108509 -480 108565 240
rect 109061 -480 109117 240
rect 109659 -480 109715 240
rect 110257 -480 110313 240
rect 110855 -480 110911 240
rect 111453 -480 111509 240
rect 112051 -480 112107 240
rect 112649 -480 112705 240
rect 113247 -480 113303 240
rect 113845 -480 113901 240
rect 114443 -480 114499 240
rect 115041 -480 115097 240
rect 115639 -480 115695 240
rect 116237 -480 116293 240
rect 116835 -480 116891 240
rect 117387 -480 117443 240
rect 117985 -480 118041 240
rect 118583 -480 118639 240
rect 119181 -480 119237 240
rect 119779 -480 119835 240
rect 120377 -480 120433 240
rect 120975 -480 121031 240
rect 121573 -480 121629 240
rect 122171 -480 122227 240
rect 122769 -480 122825 240
rect 123367 -480 123423 240
rect 123965 -480 124021 240
rect 124563 -480 124619 240
rect 125161 -480 125217 240
rect 125713 -480 125769 240
rect 126311 -480 126367 240
rect 126909 -480 126965 240
rect 127507 -480 127563 240
rect 128105 -480 128161 240
rect 128703 -480 128759 240
rect 129301 -480 129357 240
rect 129899 -480 129955 240
rect 130497 -480 130553 240
rect 131095 -480 131151 240
rect 131693 -480 131749 240
rect 132291 -480 132347 240
rect 132889 -480 132945 240
rect 133487 -480 133543 240
rect 134039 -480 134095 240
rect 134637 -480 134693 240
rect 135235 -480 135291 240
rect 135833 -480 135889 240
rect 136431 -480 136487 240
rect 137029 -480 137085 240
rect 137627 -480 137683 240
rect 138225 -480 138281 240
rect 138823 -480 138879 240
rect 139421 -480 139477 240
rect 140019 -480 140075 240
rect 140617 -480 140673 240
rect 141215 -480 141271 240
rect 141813 -480 141869 240
rect 142365 -480 142421 240
rect 142963 -480 143019 240
rect 143561 -480 143617 240
rect 144159 -480 144215 240
rect 144757 -480 144813 240
rect 145355 -480 145411 240
rect 145953 -480 146009 240
rect 146551 -480 146607 240
rect 147149 -480 147205 240
rect 147747 -480 147803 240
rect 148345 -480 148401 240
rect 148943 -480 148999 240
rect 149541 -480 149597 240
rect 150139 -480 150195 240
rect 150691 -480 150747 240
rect 151289 -480 151345 240
rect 151887 -480 151943 240
rect 152485 -480 152541 240
rect 153083 -480 153139 240
rect 153681 -480 153737 240
rect 154279 -480 154335 240
rect 154877 -480 154933 240
rect 155475 -480 155531 240
rect 156073 -480 156129 240
rect 156671 -480 156727 240
rect 157269 -480 157325 240
rect 157867 -480 157923 240
rect 158465 -480 158521 240
rect 159017 -480 159073 240
rect 159615 -480 159671 240
rect 160213 -480 160269 240
rect 160811 -480 160867 240
rect 161409 -480 161465 240
rect 162007 -480 162063 240
rect 162605 -480 162661 240
rect 163203 -480 163259 240
rect 163801 -480 163857 240
rect 164399 -480 164455 240
rect 164997 -480 165053 240
rect 165595 -480 165651 240
rect 166193 -480 166249 240
rect 166791 -480 166847 240
rect 167343 -480 167399 240
rect 167941 -480 167997 240
rect 168539 -480 168595 240
rect 169137 -480 169193 240
rect 169735 -480 169791 240
rect 170333 -480 170389 240
rect 170931 -480 170987 240
rect 171529 -480 171585 240
rect 172127 -480 172183 240
rect 172725 -480 172781 240
rect 173323 -480 173379 240
rect 173921 -480 173977 240
rect 174519 -480 174575 240
rect 175117 -480 175173 240
rect 175669 -480 175725 240
rect 176267 -480 176323 240
rect 176865 -480 176921 240
rect 177463 -480 177519 240
rect 178061 -480 178117 240
rect 178659 -480 178715 240
rect 179257 -480 179313 240
rect 179855 -480 179911 240
rect 180453 -480 180509 240
rect 181051 -480 181107 240
rect 181649 -480 181705 240
rect 182247 -480 182303 240
rect 182845 -480 182901 240
rect 183443 -480 183499 240
rect 183995 -480 184051 240
rect 184593 -480 184649 240
rect 185191 -480 185247 240
rect 185789 -480 185845 240
rect 186387 -480 186443 240
rect 186985 -480 187041 240
rect 187583 -480 187639 240
rect 188181 -480 188237 240
rect 188779 -480 188835 240
rect 189377 -480 189433 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192321 -480 192377 240
rect 192919 -480 192975 240
rect 193517 -480 193573 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197703 -480 197759 240
rect 198301 -480 198357 240
rect 198899 -480 198955 240
rect 199497 -480 199553 240
rect 200095 -480 200151 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201843 -480 201899 240
rect 202441 -480 202497 240
rect 203039 -480 203095 240
rect 203637 -480 203693 240
rect 204235 -480 204291 240
rect 204833 -480 204889 240
rect 205431 -480 205487 240
rect 206029 -480 206085 240
rect 206627 -480 206683 240
rect 207225 -480 207281 240
rect 207823 -480 207879 240
rect 208421 -480 208477 240
rect 208973 -480 209029 240
rect 209571 -480 209627 240
rect 210169 -480 210225 240
rect 210767 -480 210823 240
rect 211365 -480 211421 240
rect 211963 -480 212019 240
rect 212561 -480 212617 240
rect 213159 -480 213215 240
rect 213757 -480 213813 240
rect 214355 -480 214411 240
rect 214953 -480 215009 240
rect 215551 -480 215607 240
rect 216149 -480 216205 240
rect 216747 -480 216803 240
rect 217299 -480 217355 240
rect 217897 -480 217953 240
rect 218495 -480 218551 240
rect 219093 -480 219149 240
rect 219691 -480 219747 240
rect 220289 -480 220345 240
rect 220887 -480 220943 240
rect 221485 -480 221541 240
rect 222083 -480 222139 240
rect 222681 -480 222737 240
rect 223279 -480 223335 240
rect 223877 -480 223933 240
rect 224475 -480 224531 240
rect 225073 -480 225129 240
rect 225625 -480 225681 240
rect 226223 -480 226279 240
rect 226821 -480 226877 240
rect 227419 -480 227475 240
rect 228017 -480 228073 240
rect 228615 -480 228671 240
rect 229213 -480 229269 240
rect 229811 -480 229867 240
rect 230409 -480 230465 240
rect 231007 -480 231063 240
rect 231605 -480 231661 240
rect 232203 -480 232259 240
rect 232801 -480 232857 240
rect 233399 -480 233455 240
rect 233951 -480 234007 240
rect 234549 -480 234605 240
rect 235147 -480 235203 240
rect 235745 -480 235801 240
rect 236343 -480 236399 240
rect 236941 -480 236997 240
rect 237539 -480 237595 240
rect 238137 -480 238193 240
rect 238735 -480 238791 240
rect 239333 -480 239389 240
rect 239931 -480 239987 240
rect 240529 -480 240585 240
rect 241127 -480 241183 240
rect 241725 -480 241781 240
rect 242277 -480 242333 240
rect 242875 -480 242931 240
rect 243473 -480 243529 240
rect 244071 -480 244127 240
rect 244669 -480 244725 240
rect 245267 -480 245323 240
rect 245865 -480 245921 240
rect 246463 -480 246519 240
rect 247061 -480 247117 240
rect 247659 -480 247715 240
rect 248257 -480 248313 240
rect 248855 -480 248911 240
rect 249453 -480 249509 240
rect 250051 -480 250107 240
rect 250603 -480 250659 240
rect 251201 -480 251257 240
rect 251799 -480 251855 240
rect 252397 -480 252453 240
rect 252995 -480 253051 240
rect 253593 -480 253649 240
rect 254191 -480 254247 240
rect 254789 -480 254845 240
rect 255387 -480 255443 240
rect 255985 -480 256041 240
rect 256583 -480 256639 240
rect 257181 -480 257237 240
rect 257779 -480 257835 240
rect 258377 -480 258433 240
rect 258929 -480 258985 240
rect 259527 -480 259583 240
rect 260125 -480 260181 240
rect 260723 -480 260779 240
rect 261321 -480 261377 240
rect 261919 -480 261975 240
rect 262517 -480 262573 240
rect 263115 -480 263171 240
rect 263713 -480 263769 240
rect 264311 -480 264367 240
rect 264909 -480 264965 240
rect 265507 -480 265563 240
rect 266105 -480 266161 240
rect 266703 -480 266759 240
rect 267255 -480 267311 240
rect 267853 -480 267909 240
rect 268451 -480 268507 240
rect 269049 -480 269105 240
rect 269647 -480 269703 240
rect 270245 -480 270301 240
rect 270843 -480 270899 240
rect 271441 -480 271497 240
rect 272039 -480 272095 240
rect 272637 -480 272693 240
rect 273235 -480 273291 240
rect 273833 -480 273889 240
rect 274431 -480 274487 240
rect 275029 -480 275085 240
rect 275581 -480 275637 240
rect 276179 -480 276235 240
rect 276777 -480 276833 240
rect 277375 -480 277431 240
rect 277973 -480 278029 240
rect 278571 -480 278627 240
rect 279169 -480 279225 240
rect 279767 -480 279823 240
rect 280365 -480 280421 240
rect 280963 -480 281019 240
rect 281561 -480 281617 240
rect 282159 -480 282215 240
rect 282757 -480 282813 240
rect 283355 -480 283411 240
rect 283907 -480 283963 240
rect 284505 -480 284561 240
rect 285103 -480 285159 240
rect 285701 -480 285757 240
rect 286299 -480 286355 240
rect 286897 -480 286953 240
rect 287495 -480 287551 240
rect 288093 -480 288149 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
<<<<<<< HEAD
rect 269760 267176 270000 267236
rect 0 267040 240 267100
rect 269760 261532 270000 261592
rect 0 261192 240 261252
rect 269760 255888 270000 255948
rect 0 255344 240 255404
rect 269760 250312 270000 250372
rect 0 249428 240 249488
rect 269760 244668 270000 244728
rect 0 243580 240 243640
rect 269760 239024 270000 239084
rect 0 237732 240 237792
rect 269760 233380 270000 233440
rect 0 231816 240 231876
rect 269760 227804 270000 227864
rect 0 225968 240 226028
rect 269760 222160 270000 222220
rect 0 220120 240 220180
rect 269760 216516 270000 216576
rect 0 214204 240 214264
rect 269760 210872 270000 210932
rect 0 208356 240 208416
rect 269760 205296 270000 205356
rect 0 202508 240 202568
rect 269760 199652 270000 199712
rect 0 196592 240 196652
rect 269760 194008 270000 194068
rect 0 190744 240 190804
rect 269760 188432 270000 188492
rect 0 184896 240 184956
rect 269760 182788 270000 182848
rect 0 178980 240 179040
rect 269760 177144 270000 177204
rect 0 173132 240 173192
rect 269760 171500 270000 171560
rect 0 167284 240 167344
rect 269760 165924 270000 165984
rect 0 161368 240 161428
rect 269760 160280 270000 160340
rect 0 155520 240 155580
rect 269760 154636 270000 154696
rect 0 149672 240 149732
rect 269760 148992 270000 149052
rect 0 143756 240 143816
rect 269760 143416 270000 143476
rect 0 137908 240 137968
rect 269760 137772 270000 137832
rect 269760 132128 270000 132188
rect 0 132060 240 132120
rect 269760 126552 270000 126612
rect 0 126144 240 126204
rect 269760 120908 270000 120968
rect 0 120296 240 120356
rect 269760 115264 270000 115324
rect 0 114448 240 114508
rect 269760 109620 270000 109680
rect 0 108532 240 108592
rect 269760 104044 270000 104104
rect 0 102684 240 102744
rect 269760 98400 270000 98460
rect 0 96836 240 96896
rect 269760 92756 270000 92816
rect 0 90920 240 90980
rect 269760 87112 270000 87172
rect 0 85072 240 85132
rect 269760 81536 270000 81596
rect 0 79224 240 79284
rect 269760 75892 270000 75952
rect 0 73308 240 73368
rect 269760 70248 270000 70308
rect 0 67460 240 67520
rect 269760 64672 270000 64732
rect 0 61612 240 61672
rect 269760 59028 270000 59088
rect 0 55696 240 55756
rect 269760 53384 270000 53444
rect 0 49848 240 49908
rect 269760 47740 270000 47800
rect 0 44000 240 44060
rect 269760 42164 270000 42224
rect 0 38084 240 38144
rect 269760 36520 270000 36580
rect 0 32236 240 32296
rect 269760 30876 270000 30936
rect 0 26388 240 26448
rect 269760 25232 270000 25292
rect 0 20472 240 20532
rect 269760 19656 270000 19716
rect 0 14624 240 14684
rect 269760 14012 270000 14072
rect 0 8776 240 8836
rect 269760 8368 270000 8428
rect 0 2928 240 2988
rect 269760 2792 270000 2852
use chip-2  chip-2_0 ~/UNCCCaravel/UNCC-MPW-Shuttle/mag/tinysky
timestamp 1606345435
transform 1 0 150722 0 1 76312
box -12242 -4023 9920 9117
=======
rect 291760 348950 292480 349070
rect -480 348270 240 348390
rect 291760 343102 292480 343222
rect -480 341062 240 341182
rect 291760 337254 292480 337374
rect -480 333922 240 334042
rect 291760 331338 292480 331458
rect -480 326714 240 326834
rect 291760 325490 292480 325610
rect 291760 319642 292480 319762
rect -480 319506 240 319626
rect 291760 313794 292480 313914
rect -480 312366 240 312486
rect 291760 307878 292480 307998
rect -480 305158 240 305278
rect 291760 302030 292480 302150
rect -480 297950 240 298070
rect 291760 296182 292480 296302
rect -480 290810 240 290930
rect 291760 290334 292480 290454
rect 291760 284418 292480 284538
rect -480 283602 240 283722
rect 291760 278570 292480 278690
rect -480 276462 240 276582
rect 291760 272722 292480 272842
rect -480 269254 240 269374
rect 291760 266874 292480 266994
rect -480 262046 240 262166
rect 291760 260958 292480 261078
rect 291760 255110 292480 255230
rect -480 254906 240 255026
rect 291760 249262 292480 249382
rect -480 247698 240 247818
rect 291760 243346 292480 243466
rect -480 240490 240 240610
rect 291760 237498 292480 237618
rect -480 233350 240 233470
rect 291760 231650 292480 231770
rect -480 226142 240 226262
rect 291760 225802 292480 225922
rect 291760 219886 292480 220006
rect -480 218934 240 219054
rect 291760 214038 292480 214158
rect -480 211794 240 211914
rect 291760 208190 292480 208310
rect -480 204586 240 204706
rect 291760 202342 292480 202462
rect -480 197446 240 197566
rect 291760 196426 292480 196546
rect 291760 190578 292480 190698
rect -480 190238 240 190358
rect 291760 184730 292480 184850
rect -480 183030 240 183150
rect 291760 178882 292480 179002
rect -480 175890 240 176010
rect 291760 172966 292480 173086
rect -480 168682 240 168802
rect 291760 167118 292480 167238
rect -480 161474 240 161594
rect 291760 161270 292480 161390
rect 291760 155354 292480 155474
rect -480 154334 240 154454
rect 291760 149506 292480 149626
rect -480 147126 240 147246
rect 291760 143658 292480 143778
rect -480 139986 240 140106
rect 291760 137810 292480 137930
rect -480 132778 240 132898
rect 291760 131894 292480 132014
rect 291760 126046 292480 126166
rect -480 125570 240 125690
rect 291760 120198 292480 120318
rect -480 118430 240 118550
rect 291760 114350 292480 114470
rect -480 111222 240 111342
rect 291760 108434 292480 108554
rect -480 104014 240 104134
rect 291760 102586 292480 102706
rect -480 96874 240 96994
rect 291760 96738 292480 96858
rect 291760 90890 292480 91010
rect -480 89666 240 89786
rect 291760 84974 292480 85094
rect -480 82458 240 82578
rect 291760 79126 292480 79246
rect -480 75318 240 75438
rect 291760 73278 292480 73398
rect -480 68110 240 68230
rect 291760 67362 292480 67482
rect 291760 61514 292480 61634
rect -480 60970 240 61090
rect 291760 55666 292480 55786
rect -480 53762 240 53882
rect 291760 49818 292480 49938
rect -480 46554 240 46674
rect 291760 43902 292480 44022
rect -480 39414 240 39534
rect 291760 38054 292480 38174
rect -480 32206 240 32326
rect 291760 32206 292480 32326
rect 291760 26358 292480 26478
rect -480 24998 240 25118
rect 291760 20442 292480 20562
rect -480 17858 240 17978
rect 291760 14594 292480 14714
rect -480 10650 240 10770
rect 291760 8746 292480 8866
rect -480 3510 240 3630
rect 291760 2898 292480 3018
<< metal4 >>
rect -4218 355639 -3918 355650
rect -4218 355521 -4127 355639
rect -4009 355521 -3918 355639
rect -4218 355479 -3918 355521
rect -4218 355361 -4127 355479
rect -4009 355361 -3918 355479
rect -4218 339627 -3918 355361
rect -4218 339509 -4127 339627
rect -4009 339509 -3918 339627
rect -4218 339467 -3918 339509
rect -4218 339349 -4127 339467
rect -4009 339349 -3918 339467
rect -4218 321627 -3918 339349
rect -4218 321509 -4127 321627
rect -4009 321509 -3918 321627
rect -4218 321467 -3918 321509
rect -4218 321349 -4127 321467
rect -4009 321349 -3918 321467
rect -4218 303627 -3918 321349
rect -4218 303509 -4127 303627
rect -4009 303509 -3918 303627
rect -4218 303467 -3918 303509
rect -4218 303349 -4127 303467
rect -4009 303349 -3918 303467
rect -4218 285627 -3918 303349
rect -4218 285509 -4127 285627
rect -4009 285509 -3918 285627
rect -4218 285467 -3918 285509
rect -4218 285349 -4127 285467
rect -4009 285349 -3918 285467
rect -4218 267627 -3918 285349
rect -4218 267509 -4127 267627
rect -4009 267509 -3918 267627
rect -4218 267467 -3918 267509
rect -4218 267349 -4127 267467
rect -4009 267349 -3918 267467
rect -4218 249627 -3918 267349
rect -4218 249509 -4127 249627
rect -4009 249509 -3918 249627
rect -4218 249467 -3918 249509
rect -4218 249349 -4127 249467
rect -4009 249349 -3918 249467
rect -4218 231627 -3918 249349
rect -4218 231509 -4127 231627
rect -4009 231509 -3918 231627
rect -4218 231467 -3918 231509
rect -4218 231349 -4127 231467
rect -4009 231349 -3918 231467
rect -4218 213627 -3918 231349
rect -4218 213509 -4127 213627
rect -4009 213509 -3918 213627
rect -4218 213467 -3918 213509
rect -4218 213349 -4127 213467
rect -4009 213349 -3918 213467
rect -4218 195627 -3918 213349
rect -4218 195509 -4127 195627
rect -4009 195509 -3918 195627
rect -4218 195467 -3918 195509
rect -4218 195349 -4127 195467
rect -4009 195349 -3918 195467
rect -4218 177627 -3918 195349
rect -4218 177509 -4127 177627
rect -4009 177509 -3918 177627
rect -4218 177467 -3918 177509
rect -4218 177349 -4127 177467
rect -4009 177349 -3918 177467
rect -4218 159627 -3918 177349
rect -4218 159509 -4127 159627
rect -4009 159509 -3918 159627
rect -4218 159467 -3918 159509
rect -4218 159349 -4127 159467
rect -4009 159349 -3918 159467
rect -4218 141627 -3918 159349
rect -4218 141509 -4127 141627
rect -4009 141509 -3918 141627
rect -4218 141467 -3918 141509
rect -4218 141349 -4127 141467
rect -4009 141349 -3918 141467
rect -4218 123627 -3918 141349
rect -4218 123509 -4127 123627
rect -4009 123509 -3918 123627
rect -4218 123467 -3918 123509
rect -4218 123349 -4127 123467
rect -4009 123349 -3918 123467
rect -4218 105627 -3918 123349
rect -4218 105509 -4127 105627
rect -4009 105509 -3918 105627
rect -4218 105467 -3918 105509
rect -4218 105349 -4127 105467
rect -4009 105349 -3918 105467
rect -4218 87627 -3918 105349
rect -4218 87509 -4127 87627
rect -4009 87509 -3918 87627
rect -4218 87467 -3918 87509
rect -4218 87349 -4127 87467
rect -4009 87349 -3918 87467
rect -4218 69627 -3918 87349
rect -4218 69509 -4127 69627
rect -4009 69509 -3918 69627
rect -4218 69467 -3918 69509
rect -4218 69349 -4127 69467
rect -4009 69349 -3918 69467
rect -4218 51627 -3918 69349
rect -4218 51509 -4127 51627
rect -4009 51509 -3918 51627
rect -4218 51467 -3918 51509
rect -4218 51349 -4127 51467
rect -4009 51349 -3918 51467
rect -4218 33627 -3918 51349
rect -4218 33509 -4127 33627
rect -4009 33509 -3918 33627
rect -4218 33467 -3918 33509
rect -4218 33349 -4127 33467
rect -4009 33349 -3918 33467
rect -4218 15627 -3918 33349
rect -4218 15509 -4127 15627
rect -4009 15509 -3918 15627
rect -4218 15467 -3918 15509
rect -4218 15349 -4127 15467
rect -4009 15349 -3918 15467
rect -4218 -3393 -3918 15349
rect -3758 355179 -3458 355190
rect -3758 355061 -3667 355179
rect -3549 355061 -3458 355179
rect -3758 355019 -3458 355061
rect -3758 354901 -3667 355019
rect -3549 354901 -3458 355019
rect -3758 348627 -3458 354901
rect 5802 355179 6102 355650
rect 5802 355061 5893 355179
rect 6011 355061 6102 355179
rect 5802 355019 6102 355061
rect 5802 354901 5893 355019
rect 6011 354901 6102 355019
rect -3758 348509 -3667 348627
rect -3549 348509 -3458 348627
rect -3758 348467 -3458 348509
rect -3758 348349 -3667 348467
rect -3549 348349 -3458 348467
rect -3758 330627 -3458 348349
rect -3758 330509 -3667 330627
rect -3549 330509 -3458 330627
rect -3758 330467 -3458 330509
rect -3758 330349 -3667 330467
rect -3549 330349 -3458 330467
rect -3758 312627 -3458 330349
rect -3758 312509 -3667 312627
rect -3549 312509 -3458 312627
rect -3758 312467 -3458 312509
rect -3758 312349 -3667 312467
rect -3549 312349 -3458 312467
rect -3758 294627 -3458 312349
rect -3758 294509 -3667 294627
rect -3549 294509 -3458 294627
rect -3758 294467 -3458 294509
rect -3758 294349 -3667 294467
rect -3549 294349 -3458 294467
rect -3758 276627 -3458 294349
rect -3758 276509 -3667 276627
rect -3549 276509 -3458 276627
rect -3758 276467 -3458 276509
rect -3758 276349 -3667 276467
rect -3549 276349 -3458 276467
rect -3758 258627 -3458 276349
rect -3758 258509 -3667 258627
rect -3549 258509 -3458 258627
rect -3758 258467 -3458 258509
rect -3758 258349 -3667 258467
rect -3549 258349 -3458 258467
rect -3758 240627 -3458 258349
rect -3758 240509 -3667 240627
rect -3549 240509 -3458 240627
rect -3758 240467 -3458 240509
rect -3758 240349 -3667 240467
rect -3549 240349 -3458 240467
rect -3758 222627 -3458 240349
rect -3758 222509 -3667 222627
rect -3549 222509 -3458 222627
rect -3758 222467 -3458 222509
rect -3758 222349 -3667 222467
rect -3549 222349 -3458 222467
rect -3758 204627 -3458 222349
rect -3758 204509 -3667 204627
rect -3549 204509 -3458 204627
rect -3758 204467 -3458 204509
rect -3758 204349 -3667 204467
rect -3549 204349 -3458 204467
rect -3758 186627 -3458 204349
rect -3758 186509 -3667 186627
rect -3549 186509 -3458 186627
rect -3758 186467 -3458 186509
rect -3758 186349 -3667 186467
rect -3549 186349 -3458 186467
rect -3758 168627 -3458 186349
rect -3758 168509 -3667 168627
rect -3549 168509 -3458 168627
rect -3758 168467 -3458 168509
rect -3758 168349 -3667 168467
rect -3549 168349 -3458 168467
rect -3758 150627 -3458 168349
rect -3758 150509 -3667 150627
rect -3549 150509 -3458 150627
rect -3758 150467 -3458 150509
rect -3758 150349 -3667 150467
rect -3549 150349 -3458 150467
rect -3758 132627 -3458 150349
rect -3758 132509 -3667 132627
rect -3549 132509 -3458 132627
rect -3758 132467 -3458 132509
rect -3758 132349 -3667 132467
rect -3549 132349 -3458 132467
rect -3758 114627 -3458 132349
rect -3758 114509 -3667 114627
rect -3549 114509 -3458 114627
rect -3758 114467 -3458 114509
rect -3758 114349 -3667 114467
rect -3549 114349 -3458 114467
rect -3758 96627 -3458 114349
rect -3758 96509 -3667 96627
rect -3549 96509 -3458 96627
rect -3758 96467 -3458 96509
rect -3758 96349 -3667 96467
rect -3549 96349 -3458 96467
rect -3758 78627 -3458 96349
rect -3758 78509 -3667 78627
rect -3549 78509 -3458 78627
rect -3758 78467 -3458 78509
rect -3758 78349 -3667 78467
rect -3549 78349 -3458 78467
rect -3758 60627 -3458 78349
rect -3758 60509 -3667 60627
rect -3549 60509 -3458 60627
rect -3758 60467 -3458 60509
rect -3758 60349 -3667 60467
rect -3549 60349 -3458 60467
rect -3758 42627 -3458 60349
rect -3758 42509 -3667 42627
rect -3549 42509 -3458 42627
rect -3758 42467 -3458 42509
rect -3758 42349 -3667 42467
rect -3549 42349 -3458 42467
rect -3758 24627 -3458 42349
rect -3758 24509 -3667 24627
rect -3549 24509 -3458 24627
rect -3758 24467 -3458 24509
rect -3758 24349 -3667 24467
rect -3549 24349 -3458 24467
rect -3758 6627 -3458 24349
rect -3758 6509 -3667 6627
rect -3549 6509 -3458 6627
rect -3758 6467 -3458 6509
rect -3758 6349 -3667 6467
rect -3549 6349 -3458 6467
rect -3758 -2933 -3458 6349
rect -3298 354719 -2998 354730
rect -3298 354601 -3207 354719
rect -3089 354601 -2998 354719
rect -3298 354559 -2998 354601
rect -3298 354441 -3207 354559
rect -3089 354441 -2998 354559
rect -3298 337827 -2998 354441
rect -3298 337709 -3207 337827
rect -3089 337709 -2998 337827
rect -3298 337667 -2998 337709
rect -3298 337549 -3207 337667
rect -3089 337549 -2998 337667
rect -3298 319827 -2998 337549
rect -3298 319709 -3207 319827
rect -3089 319709 -2998 319827
rect -3298 319667 -2998 319709
rect -3298 319549 -3207 319667
rect -3089 319549 -2998 319667
rect -3298 301827 -2998 319549
rect -3298 301709 -3207 301827
rect -3089 301709 -2998 301827
rect -3298 301667 -2998 301709
rect -3298 301549 -3207 301667
rect -3089 301549 -2998 301667
rect -3298 283827 -2998 301549
rect -3298 283709 -3207 283827
rect -3089 283709 -2998 283827
rect -3298 283667 -2998 283709
rect -3298 283549 -3207 283667
rect -3089 283549 -2998 283667
rect -3298 265827 -2998 283549
rect -3298 265709 -3207 265827
rect -3089 265709 -2998 265827
rect -3298 265667 -2998 265709
rect -3298 265549 -3207 265667
rect -3089 265549 -2998 265667
rect -3298 247827 -2998 265549
rect -3298 247709 -3207 247827
rect -3089 247709 -2998 247827
rect -3298 247667 -2998 247709
rect -3298 247549 -3207 247667
rect -3089 247549 -2998 247667
rect -3298 229827 -2998 247549
rect -3298 229709 -3207 229827
rect -3089 229709 -2998 229827
rect -3298 229667 -2998 229709
rect -3298 229549 -3207 229667
rect -3089 229549 -2998 229667
rect -3298 211827 -2998 229549
rect -3298 211709 -3207 211827
rect -3089 211709 -2998 211827
rect -3298 211667 -2998 211709
rect -3298 211549 -3207 211667
rect -3089 211549 -2998 211667
rect -3298 193827 -2998 211549
rect -3298 193709 -3207 193827
rect -3089 193709 -2998 193827
rect -3298 193667 -2998 193709
rect -3298 193549 -3207 193667
rect -3089 193549 -2998 193667
rect -3298 175827 -2998 193549
rect -3298 175709 -3207 175827
rect -3089 175709 -2998 175827
rect -3298 175667 -2998 175709
rect -3298 175549 -3207 175667
rect -3089 175549 -2998 175667
rect -3298 157827 -2998 175549
rect -3298 157709 -3207 157827
rect -3089 157709 -2998 157827
rect -3298 157667 -2998 157709
rect -3298 157549 -3207 157667
rect -3089 157549 -2998 157667
rect -3298 139827 -2998 157549
rect -3298 139709 -3207 139827
rect -3089 139709 -2998 139827
rect -3298 139667 -2998 139709
rect -3298 139549 -3207 139667
rect -3089 139549 -2998 139667
rect -3298 121827 -2998 139549
rect -3298 121709 -3207 121827
rect -3089 121709 -2998 121827
rect -3298 121667 -2998 121709
rect -3298 121549 -3207 121667
rect -3089 121549 -2998 121667
rect -3298 103827 -2998 121549
rect -3298 103709 -3207 103827
rect -3089 103709 -2998 103827
rect -3298 103667 -2998 103709
rect -3298 103549 -3207 103667
rect -3089 103549 -2998 103667
rect -3298 85827 -2998 103549
rect -3298 85709 -3207 85827
rect -3089 85709 -2998 85827
rect -3298 85667 -2998 85709
rect -3298 85549 -3207 85667
rect -3089 85549 -2998 85667
rect -3298 67827 -2998 85549
rect -3298 67709 -3207 67827
rect -3089 67709 -2998 67827
rect -3298 67667 -2998 67709
rect -3298 67549 -3207 67667
rect -3089 67549 -2998 67667
rect -3298 49827 -2998 67549
rect -3298 49709 -3207 49827
rect -3089 49709 -2998 49827
rect -3298 49667 -2998 49709
rect -3298 49549 -3207 49667
rect -3089 49549 -2998 49667
rect -3298 31827 -2998 49549
rect -3298 31709 -3207 31827
rect -3089 31709 -2998 31827
rect -3298 31667 -2998 31709
rect -3298 31549 -3207 31667
rect -3089 31549 -2998 31667
rect -3298 13827 -2998 31549
rect -3298 13709 -3207 13827
rect -3089 13709 -2998 13827
rect -3298 13667 -2998 13709
rect -3298 13549 -3207 13667
rect -3089 13549 -2998 13667
rect -3298 -2473 -2998 13549
rect -2838 354259 -2538 354270
rect -2838 354141 -2747 354259
rect -2629 354141 -2538 354259
rect -2838 354099 -2538 354141
rect -2838 353981 -2747 354099
rect -2629 353981 -2538 354099
rect -2838 346827 -2538 353981
rect 4002 354259 4302 354730
rect 4002 354141 4093 354259
rect 4211 354141 4302 354259
rect 4002 354099 4302 354141
rect 4002 353981 4093 354099
rect 4211 353981 4302 354099
rect -2838 346709 -2747 346827
rect -2629 346709 -2538 346827
rect -2838 346667 -2538 346709
rect -2838 346549 -2747 346667
rect -2629 346549 -2538 346667
rect -2838 328827 -2538 346549
rect -2838 328709 -2747 328827
rect -2629 328709 -2538 328827
rect -2838 328667 -2538 328709
rect -2838 328549 -2747 328667
rect -2629 328549 -2538 328667
rect -2838 310827 -2538 328549
rect -2838 310709 -2747 310827
rect -2629 310709 -2538 310827
rect -2838 310667 -2538 310709
rect -2838 310549 -2747 310667
rect -2629 310549 -2538 310667
rect -2838 292827 -2538 310549
rect -2838 292709 -2747 292827
rect -2629 292709 -2538 292827
rect -2838 292667 -2538 292709
rect -2838 292549 -2747 292667
rect -2629 292549 -2538 292667
rect -2838 274827 -2538 292549
rect -2838 274709 -2747 274827
rect -2629 274709 -2538 274827
rect -2838 274667 -2538 274709
rect -2838 274549 -2747 274667
rect -2629 274549 -2538 274667
rect -2838 256827 -2538 274549
rect -2838 256709 -2747 256827
rect -2629 256709 -2538 256827
rect -2838 256667 -2538 256709
rect -2838 256549 -2747 256667
rect -2629 256549 -2538 256667
rect -2838 238827 -2538 256549
rect -2838 238709 -2747 238827
rect -2629 238709 -2538 238827
rect -2838 238667 -2538 238709
rect -2838 238549 -2747 238667
rect -2629 238549 -2538 238667
rect -2838 220827 -2538 238549
rect -2838 220709 -2747 220827
rect -2629 220709 -2538 220827
rect -2838 220667 -2538 220709
rect -2838 220549 -2747 220667
rect -2629 220549 -2538 220667
rect -2838 202827 -2538 220549
rect -2838 202709 -2747 202827
rect -2629 202709 -2538 202827
rect -2838 202667 -2538 202709
rect -2838 202549 -2747 202667
rect -2629 202549 -2538 202667
rect -2838 184827 -2538 202549
rect -2838 184709 -2747 184827
rect -2629 184709 -2538 184827
rect -2838 184667 -2538 184709
rect -2838 184549 -2747 184667
rect -2629 184549 -2538 184667
rect -2838 166827 -2538 184549
rect -2838 166709 -2747 166827
rect -2629 166709 -2538 166827
rect -2838 166667 -2538 166709
rect -2838 166549 -2747 166667
rect -2629 166549 -2538 166667
rect -2838 148827 -2538 166549
rect -2838 148709 -2747 148827
rect -2629 148709 -2538 148827
rect -2838 148667 -2538 148709
rect -2838 148549 -2747 148667
rect -2629 148549 -2538 148667
rect -2838 130827 -2538 148549
rect -2838 130709 -2747 130827
rect -2629 130709 -2538 130827
rect -2838 130667 -2538 130709
rect -2838 130549 -2747 130667
rect -2629 130549 -2538 130667
rect -2838 112827 -2538 130549
rect -2838 112709 -2747 112827
rect -2629 112709 -2538 112827
rect -2838 112667 -2538 112709
rect -2838 112549 -2747 112667
rect -2629 112549 -2538 112667
rect -2838 94827 -2538 112549
rect -2838 94709 -2747 94827
rect -2629 94709 -2538 94827
rect -2838 94667 -2538 94709
rect -2838 94549 -2747 94667
rect -2629 94549 -2538 94667
rect -2838 76827 -2538 94549
rect -2838 76709 -2747 76827
rect -2629 76709 -2538 76827
rect -2838 76667 -2538 76709
rect -2838 76549 -2747 76667
rect -2629 76549 -2538 76667
rect -2838 58827 -2538 76549
rect -2838 58709 -2747 58827
rect -2629 58709 -2538 58827
rect -2838 58667 -2538 58709
rect -2838 58549 -2747 58667
rect -2629 58549 -2538 58667
rect -2838 40827 -2538 58549
rect -2838 40709 -2747 40827
rect -2629 40709 -2538 40827
rect -2838 40667 -2538 40709
rect -2838 40549 -2747 40667
rect -2629 40549 -2538 40667
rect -2838 22827 -2538 40549
rect -2838 22709 -2747 22827
rect -2629 22709 -2538 22827
rect -2838 22667 -2538 22709
rect -2838 22549 -2747 22667
rect -2629 22549 -2538 22667
rect -2838 4827 -2538 22549
rect -2838 4709 -2747 4827
rect -2629 4709 -2538 4827
rect -2838 4667 -2538 4709
rect -2838 4549 -2747 4667
rect -2629 4549 -2538 4667
rect -2838 -2013 -2538 4549
rect -2378 353799 -2078 353810
rect -2378 353681 -2287 353799
rect -2169 353681 -2078 353799
rect -2378 353639 -2078 353681
rect -2378 353521 -2287 353639
rect -2169 353521 -2078 353639
rect -2378 336027 -2078 353521
rect -2378 335909 -2287 336027
rect -2169 335909 -2078 336027
rect -2378 335867 -2078 335909
rect -2378 335749 -2287 335867
rect -2169 335749 -2078 335867
rect -2378 318027 -2078 335749
rect -2378 317909 -2287 318027
rect -2169 317909 -2078 318027
rect -2378 317867 -2078 317909
rect -2378 317749 -2287 317867
rect -2169 317749 -2078 317867
rect -2378 300027 -2078 317749
rect -2378 299909 -2287 300027
rect -2169 299909 -2078 300027
rect -2378 299867 -2078 299909
rect -2378 299749 -2287 299867
rect -2169 299749 -2078 299867
rect -2378 282027 -2078 299749
rect -2378 281909 -2287 282027
rect -2169 281909 -2078 282027
rect -2378 281867 -2078 281909
rect -2378 281749 -2287 281867
rect -2169 281749 -2078 281867
rect -2378 264027 -2078 281749
rect -2378 263909 -2287 264027
rect -2169 263909 -2078 264027
rect -2378 263867 -2078 263909
rect -2378 263749 -2287 263867
rect -2169 263749 -2078 263867
rect -2378 246027 -2078 263749
rect -2378 245909 -2287 246027
rect -2169 245909 -2078 246027
rect -2378 245867 -2078 245909
rect -2378 245749 -2287 245867
rect -2169 245749 -2078 245867
rect -2378 228027 -2078 245749
rect -2378 227909 -2287 228027
rect -2169 227909 -2078 228027
rect -2378 227867 -2078 227909
rect -2378 227749 -2287 227867
rect -2169 227749 -2078 227867
rect -2378 210027 -2078 227749
rect -2378 209909 -2287 210027
rect -2169 209909 -2078 210027
rect -2378 209867 -2078 209909
rect -2378 209749 -2287 209867
rect -2169 209749 -2078 209867
rect -2378 192027 -2078 209749
rect -2378 191909 -2287 192027
rect -2169 191909 -2078 192027
rect -2378 191867 -2078 191909
rect -2378 191749 -2287 191867
rect -2169 191749 -2078 191867
rect -2378 174027 -2078 191749
rect -2378 173909 -2287 174027
rect -2169 173909 -2078 174027
rect -2378 173867 -2078 173909
rect -2378 173749 -2287 173867
rect -2169 173749 -2078 173867
rect -2378 156027 -2078 173749
rect -2378 155909 -2287 156027
rect -2169 155909 -2078 156027
rect -2378 155867 -2078 155909
rect -2378 155749 -2287 155867
rect -2169 155749 -2078 155867
rect -2378 138027 -2078 155749
rect -2378 137909 -2287 138027
rect -2169 137909 -2078 138027
rect -2378 137867 -2078 137909
rect -2378 137749 -2287 137867
rect -2169 137749 -2078 137867
rect -2378 120027 -2078 137749
rect -2378 119909 -2287 120027
rect -2169 119909 -2078 120027
rect -2378 119867 -2078 119909
rect -2378 119749 -2287 119867
rect -2169 119749 -2078 119867
rect -2378 102027 -2078 119749
rect -2378 101909 -2287 102027
rect -2169 101909 -2078 102027
rect -2378 101867 -2078 101909
rect -2378 101749 -2287 101867
rect -2169 101749 -2078 101867
rect -2378 84027 -2078 101749
rect -2378 83909 -2287 84027
rect -2169 83909 -2078 84027
rect -2378 83867 -2078 83909
rect -2378 83749 -2287 83867
rect -2169 83749 -2078 83867
rect -2378 66027 -2078 83749
rect -2378 65909 -2287 66027
rect -2169 65909 -2078 66027
rect -2378 65867 -2078 65909
rect -2378 65749 -2287 65867
rect -2169 65749 -2078 65867
rect -2378 48027 -2078 65749
rect -2378 47909 -2287 48027
rect -2169 47909 -2078 48027
rect -2378 47867 -2078 47909
rect -2378 47749 -2287 47867
rect -2169 47749 -2078 47867
rect -2378 30027 -2078 47749
rect -2378 29909 -2287 30027
rect -2169 29909 -2078 30027
rect -2378 29867 -2078 29909
rect -2378 29749 -2287 29867
rect -2169 29749 -2078 29867
rect -2378 12027 -2078 29749
rect -2378 11909 -2287 12027
rect -2169 11909 -2078 12027
rect -2378 11867 -2078 11909
rect -2378 11749 -2287 11867
rect -2169 11749 -2078 11867
rect -2378 -1553 -2078 11749
rect -1918 353339 -1618 353350
rect -1918 353221 -1827 353339
rect -1709 353221 -1618 353339
rect -1918 353179 -1618 353221
rect -1918 353061 -1827 353179
rect -1709 353061 -1618 353179
rect -1918 345027 -1618 353061
rect 2202 353339 2502 353810
rect 2202 353221 2293 353339
rect 2411 353221 2502 353339
rect 2202 353179 2502 353221
rect 2202 353061 2293 353179
rect 2411 353061 2502 353179
rect -1918 344909 -1827 345027
rect -1709 344909 -1618 345027
rect -1918 344867 -1618 344909
rect -1918 344749 -1827 344867
rect -1709 344749 -1618 344867
rect -1918 327027 -1618 344749
rect -1918 326909 -1827 327027
rect -1709 326909 -1618 327027
rect -1918 326867 -1618 326909
rect -1918 326749 -1827 326867
rect -1709 326749 -1618 326867
rect -1918 309027 -1618 326749
rect -1918 308909 -1827 309027
rect -1709 308909 -1618 309027
rect -1918 308867 -1618 308909
rect -1918 308749 -1827 308867
rect -1709 308749 -1618 308867
rect -1918 291027 -1618 308749
rect -1918 290909 -1827 291027
rect -1709 290909 -1618 291027
rect -1918 290867 -1618 290909
rect -1918 290749 -1827 290867
rect -1709 290749 -1618 290867
rect -1918 273027 -1618 290749
rect -1918 272909 -1827 273027
rect -1709 272909 -1618 273027
rect -1918 272867 -1618 272909
rect -1918 272749 -1827 272867
rect -1709 272749 -1618 272867
rect -1918 255027 -1618 272749
rect -1918 254909 -1827 255027
rect -1709 254909 -1618 255027
rect -1918 254867 -1618 254909
rect -1918 254749 -1827 254867
rect -1709 254749 -1618 254867
rect -1918 237027 -1618 254749
rect -1918 236909 -1827 237027
rect -1709 236909 -1618 237027
rect -1918 236867 -1618 236909
rect -1918 236749 -1827 236867
rect -1709 236749 -1618 236867
rect -1918 219027 -1618 236749
rect -1918 218909 -1827 219027
rect -1709 218909 -1618 219027
rect -1918 218867 -1618 218909
rect -1918 218749 -1827 218867
rect -1709 218749 -1618 218867
rect -1918 201027 -1618 218749
rect -1918 200909 -1827 201027
rect -1709 200909 -1618 201027
rect -1918 200867 -1618 200909
rect -1918 200749 -1827 200867
rect -1709 200749 -1618 200867
rect -1918 183027 -1618 200749
rect -1918 182909 -1827 183027
rect -1709 182909 -1618 183027
rect -1918 182867 -1618 182909
rect -1918 182749 -1827 182867
rect -1709 182749 -1618 182867
rect -1918 165027 -1618 182749
rect -1918 164909 -1827 165027
rect -1709 164909 -1618 165027
rect -1918 164867 -1618 164909
rect -1918 164749 -1827 164867
rect -1709 164749 -1618 164867
rect -1918 147027 -1618 164749
rect -1918 146909 -1827 147027
rect -1709 146909 -1618 147027
rect -1918 146867 -1618 146909
rect -1918 146749 -1827 146867
rect -1709 146749 -1618 146867
rect -1918 129027 -1618 146749
rect -1918 128909 -1827 129027
rect -1709 128909 -1618 129027
rect -1918 128867 -1618 128909
rect -1918 128749 -1827 128867
rect -1709 128749 -1618 128867
rect -1918 111027 -1618 128749
rect -1918 110909 -1827 111027
rect -1709 110909 -1618 111027
rect -1918 110867 -1618 110909
rect -1918 110749 -1827 110867
rect -1709 110749 -1618 110867
rect -1918 93027 -1618 110749
rect -1918 92909 -1827 93027
rect -1709 92909 -1618 93027
rect -1918 92867 -1618 92909
rect -1918 92749 -1827 92867
rect -1709 92749 -1618 92867
rect -1918 75027 -1618 92749
rect -1918 74909 -1827 75027
rect -1709 74909 -1618 75027
rect -1918 74867 -1618 74909
rect -1918 74749 -1827 74867
rect -1709 74749 -1618 74867
rect -1918 57027 -1618 74749
rect -1918 56909 -1827 57027
rect -1709 56909 -1618 57027
rect -1918 56867 -1618 56909
rect -1918 56749 -1827 56867
rect -1709 56749 -1618 56867
rect -1918 39027 -1618 56749
rect -1918 38909 -1827 39027
rect -1709 38909 -1618 39027
rect -1918 38867 -1618 38909
rect -1918 38749 -1827 38867
rect -1709 38749 -1618 38867
rect -1918 21027 -1618 38749
rect -1918 20909 -1827 21027
rect -1709 20909 -1618 21027
rect -1918 20867 -1618 20909
rect -1918 20749 -1827 20867
rect -1709 20749 -1618 20867
rect -1918 3027 -1618 20749
rect -1918 2909 -1827 3027
rect -1709 2909 -1618 3027
rect -1918 2867 -1618 2909
rect -1918 2749 -1827 2867
rect -1709 2749 -1618 2867
rect -1918 -1093 -1618 2749
rect -1458 352879 -1158 352890
rect -1458 352761 -1367 352879
rect -1249 352761 -1158 352879
rect -1458 352719 -1158 352761
rect -1458 352601 -1367 352719
rect -1249 352601 -1158 352719
rect -1458 334227 -1158 352601
rect -1458 334109 -1367 334227
rect -1249 334109 -1158 334227
rect -1458 334067 -1158 334109
rect -1458 333949 -1367 334067
rect -1249 333949 -1158 334067
rect -1458 316227 -1158 333949
rect -1458 316109 -1367 316227
rect -1249 316109 -1158 316227
rect -1458 316067 -1158 316109
rect -1458 315949 -1367 316067
rect -1249 315949 -1158 316067
rect -1458 298227 -1158 315949
rect -1458 298109 -1367 298227
rect -1249 298109 -1158 298227
rect -1458 298067 -1158 298109
rect -1458 297949 -1367 298067
rect -1249 297949 -1158 298067
rect -1458 280227 -1158 297949
rect -1458 280109 -1367 280227
rect -1249 280109 -1158 280227
rect -1458 280067 -1158 280109
rect -1458 279949 -1367 280067
rect -1249 279949 -1158 280067
rect -1458 262227 -1158 279949
rect -1458 262109 -1367 262227
rect -1249 262109 -1158 262227
rect -1458 262067 -1158 262109
rect -1458 261949 -1367 262067
rect -1249 261949 -1158 262067
rect -1458 244227 -1158 261949
rect -1458 244109 -1367 244227
rect -1249 244109 -1158 244227
rect -1458 244067 -1158 244109
rect -1458 243949 -1367 244067
rect -1249 243949 -1158 244067
rect -1458 226227 -1158 243949
rect -1458 226109 -1367 226227
rect -1249 226109 -1158 226227
rect -1458 226067 -1158 226109
rect -1458 225949 -1367 226067
rect -1249 225949 -1158 226067
rect -1458 208227 -1158 225949
rect -1458 208109 -1367 208227
rect -1249 208109 -1158 208227
rect -1458 208067 -1158 208109
rect -1458 207949 -1367 208067
rect -1249 207949 -1158 208067
rect -1458 190227 -1158 207949
rect -1458 190109 -1367 190227
rect -1249 190109 -1158 190227
rect -1458 190067 -1158 190109
rect -1458 189949 -1367 190067
rect -1249 189949 -1158 190067
rect -1458 172227 -1158 189949
rect -1458 172109 -1367 172227
rect -1249 172109 -1158 172227
rect -1458 172067 -1158 172109
rect -1458 171949 -1367 172067
rect -1249 171949 -1158 172067
rect -1458 154227 -1158 171949
rect -1458 154109 -1367 154227
rect -1249 154109 -1158 154227
rect -1458 154067 -1158 154109
rect -1458 153949 -1367 154067
rect -1249 153949 -1158 154067
rect -1458 136227 -1158 153949
rect -1458 136109 -1367 136227
rect -1249 136109 -1158 136227
rect -1458 136067 -1158 136109
rect -1458 135949 -1367 136067
rect -1249 135949 -1158 136067
rect -1458 118227 -1158 135949
rect -1458 118109 -1367 118227
rect -1249 118109 -1158 118227
rect -1458 118067 -1158 118109
rect -1458 117949 -1367 118067
rect -1249 117949 -1158 118067
rect -1458 100227 -1158 117949
rect -1458 100109 -1367 100227
rect -1249 100109 -1158 100227
rect -1458 100067 -1158 100109
rect -1458 99949 -1367 100067
rect -1249 99949 -1158 100067
rect -1458 82227 -1158 99949
rect -1458 82109 -1367 82227
rect -1249 82109 -1158 82227
rect -1458 82067 -1158 82109
rect -1458 81949 -1367 82067
rect -1249 81949 -1158 82067
rect -1458 64227 -1158 81949
rect -1458 64109 -1367 64227
rect -1249 64109 -1158 64227
rect -1458 64067 -1158 64109
rect -1458 63949 -1367 64067
rect -1249 63949 -1158 64067
rect -1458 46227 -1158 63949
rect -1458 46109 -1367 46227
rect -1249 46109 -1158 46227
rect -1458 46067 -1158 46109
rect -1458 45949 -1367 46067
rect -1249 45949 -1158 46067
rect -1458 28227 -1158 45949
rect -1458 28109 -1367 28227
rect -1249 28109 -1158 28227
rect -1458 28067 -1158 28109
rect -1458 27949 -1367 28067
rect -1249 27949 -1158 28067
rect -1458 10227 -1158 27949
rect -1458 10109 -1367 10227
rect -1249 10109 -1158 10227
rect -1458 10067 -1158 10109
rect -1458 9949 -1367 10067
rect -1249 9949 -1158 10067
rect -1458 -633 -1158 9949
rect -998 352419 -698 352430
rect -998 352301 -907 352419
rect -789 352301 -698 352419
rect -998 352259 -698 352301
rect -998 352141 -907 352259
rect -789 352141 -698 352259
rect -998 343227 -698 352141
rect 402 352419 702 352890
rect 402 352301 493 352419
rect 611 352301 702 352419
rect 402 352259 702 352301
rect 402 352141 493 352259
rect 611 352141 702 352259
rect 402 351760 702 352141
rect 2202 351760 2502 353061
rect 4002 351760 4302 353981
rect 5802 351760 6102 354901
rect 14802 355639 15102 355650
rect 14802 355521 14893 355639
rect 15011 355521 15102 355639
rect 14802 355479 15102 355521
rect 14802 355361 14893 355479
rect 15011 355361 15102 355479
rect 13002 354719 13302 354730
rect 13002 354601 13093 354719
rect 13211 354601 13302 354719
rect 13002 354559 13302 354601
rect 13002 354441 13093 354559
rect 13211 354441 13302 354559
rect 11202 353799 11502 353810
rect 11202 353681 11293 353799
rect 11411 353681 11502 353799
rect 11202 353639 11502 353681
rect 11202 353521 11293 353639
rect 11411 353521 11502 353639
rect 9402 352879 9702 352890
rect 9402 352761 9493 352879
rect 9611 352761 9702 352879
rect 9402 352719 9702 352761
rect 9402 352601 9493 352719
rect 9611 352601 9702 352719
rect 9402 351760 9702 352601
rect 11202 351760 11502 353521
rect 13002 351760 13302 354441
rect 14802 351760 15102 355361
rect 23802 355179 24102 355650
rect 23802 355061 23893 355179
rect 24011 355061 24102 355179
rect 23802 355019 24102 355061
rect 23802 354901 23893 355019
rect 24011 354901 24102 355019
rect 22002 354259 22302 354730
rect 22002 354141 22093 354259
rect 22211 354141 22302 354259
rect 22002 354099 22302 354141
rect 22002 353981 22093 354099
rect 22211 353981 22302 354099
rect 20202 353339 20502 353810
rect 20202 353221 20293 353339
rect 20411 353221 20502 353339
rect 20202 353179 20502 353221
rect 20202 353061 20293 353179
rect 20411 353061 20502 353179
rect 18402 352419 18702 352890
rect 18402 352301 18493 352419
rect 18611 352301 18702 352419
rect 18402 352259 18702 352301
rect 18402 352141 18493 352259
rect 18611 352141 18702 352259
rect 18402 351760 18702 352141
rect 20202 351760 20502 353061
rect 22002 351760 22302 353981
rect 23802 351760 24102 354901
rect 32802 355639 33102 355650
rect 32802 355521 32893 355639
rect 33011 355521 33102 355639
rect 32802 355479 33102 355521
rect 32802 355361 32893 355479
rect 33011 355361 33102 355479
rect 31002 354719 31302 354730
rect 31002 354601 31093 354719
rect 31211 354601 31302 354719
rect 31002 354559 31302 354601
rect 31002 354441 31093 354559
rect 31211 354441 31302 354559
rect 29202 353799 29502 353810
rect 29202 353681 29293 353799
rect 29411 353681 29502 353799
rect 29202 353639 29502 353681
rect 29202 353521 29293 353639
rect 29411 353521 29502 353639
rect 27402 352879 27702 352890
rect 27402 352761 27493 352879
rect 27611 352761 27702 352879
rect 27402 352719 27702 352761
rect 27402 352601 27493 352719
rect 27611 352601 27702 352719
rect 27402 351760 27702 352601
rect 29202 351760 29502 353521
rect 31002 351760 31302 354441
rect 32802 351760 33102 355361
rect 41802 355179 42102 355650
rect 41802 355061 41893 355179
rect 42011 355061 42102 355179
rect 41802 355019 42102 355061
rect 41802 354901 41893 355019
rect 42011 354901 42102 355019
rect 40002 354259 40302 354730
rect 40002 354141 40093 354259
rect 40211 354141 40302 354259
rect 40002 354099 40302 354141
rect 40002 353981 40093 354099
rect 40211 353981 40302 354099
rect 38202 353339 38502 353810
rect 38202 353221 38293 353339
rect 38411 353221 38502 353339
rect 38202 353179 38502 353221
rect 38202 353061 38293 353179
rect 38411 353061 38502 353179
rect 36402 352419 36702 352890
rect 36402 352301 36493 352419
rect 36611 352301 36702 352419
rect 36402 352259 36702 352301
rect 36402 352141 36493 352259
rect 36611 352141 36702 352259
rect 36402 351760 36702 352141
rect 38202 351760 38502 353061
rect 40002 351760 40302 353981
rect 41802 351760 42102 354901
rect 50802 355639 51102 355650
rect 50802 355521 50893 355639
rect 51011 355521 51102 355639
rect 50802 355479 51102 355521
rect 50802 355361 50893 355479
rect 51011 355361 51102 355479
rect 49002 354719 49302 354730
rect 49002 354601 49093 354719
rect 49211 354601 49302 354719
rect 49002 354559 49302 354601
rect 49002 354441 49093 354559
rect 49211 354441 49302 354559
rect 47202 353799 47502 353810
rect 47202 353681 47293 353799
rect 47411 353681 47502 353799
rect 47202 353639 47502 353681
rect 47202 353521 47293 353639
rect 47411 353521 47502 353639
rect 45402 352879 45702 352890
rect 45402 352761 45493 352879
rect 45611 352761 45702 352879
rect 45402 352719 45702 352761
rect 45402 352601 45493 352719
rect 45611 352601 45702 352719
rect 45402 351760 45702 352601
rect 47202 351760 47502 353521
rect 49002 351760 49302 354441
rect 50802 351760 51102 355361
rect 59802 355179 60102 355650
rect 59802 355061 59893 355179
rect 60011 355061 60102 355179
rect 59802 355019 60102 355061
rect 59802 354901 59893 355019
rect 60011 354901 60102 355019
rect 58002 354259 58302 354730
rect 58002 354141 58093 354259
rect 58211 354141 58302 354259
rect 58002 354099 58302 354141
rect 58002 353981 58093 354099
rect 58211 353981 58302 354099
rect 56202 353339 56502 353810
rect 56202 353221 56293 353339
rect 56411 353221 56502 353339
rect 56202 353179 56502 353221
rect 56202 353061 56293 353179
rect 56411 353061 56502 353179
rect 54402 352419 54702 352890
rect 54402 352301 54493 352419
rect 54611 352301 54702 352419
rect 54402 352259 54702 352301
rect 54402 352141 54493 352259
rect 54611 352141 54702 352259
rect 54402 351760 54702 352141
rect 56202 351760 56502 353061
rect 58002 351760 58302 353981
rect 59802 351760 60102 354901
rect 68802 355639 69102 355650
rect 68802 355521 68893 355639
rect 69011 355521 69102 355639
rect 68802 355479 69102 355521
rect 68802 355361 68893 355479
rect 69011 355361 69102 355479
rect 67002 354719 67302 354730
rect 67002 354601 67093 354719
rect 67211 354601 67302 354719
rect 67002 354559 67302 354601
rect 67002 354441 67093 354559
rect 67211 354441 67302 354559
rect 65202 353799 65502 353810
rect 65202 353681 65293 353799
rect 65411 353681 65502 353799
rect 65202 353639 65502 353681
rect 65202 353521 65293 353639
rect 65411 353521 65502 353639
rect 63402 352879 63702 352890
rect 63402 352761 63493 352879
rect 63611 352761 63702 352879
rect 63402 352719 63702 352761
rect 63402 352601 63493 352719
rect 63611 352601 63702 352719
rect 63402 351760 63702 352601
rect 65202 351760 65502 353521
rect 67002 351760 67302 354441
rect 68802 351760 69102 355361
rect 77802 355179 78102 355650
rect 77802 355061 77893 355179
rect 78011 355061 78102 355179
rect 77802 355019 78102 355061
rect 77802 354901 77893 355019
rect 78011 354901 78102 355019
rect 76002 354259 76302 354730
rect 76002 354141 76093 354259
rect 76211 354141 76302 354259
rect 76002 354099 76302 354141
rect 76002 353981 76093 354099
rect 76211 353981 76302 354099
rect 74202 353339 74502 353810
rect 74202 353221 74293 353339
rect 74411 353221 74502 353339
rect 74202 353179 74502 353221
rect 74202 353061 74293 353179
rect 74411 353061 74502 353179
rect 72402 352419 72702 352890
rect 72402 352301 72493 352419
rect 72611 352301 72702 352419
rect 72402 352259 72702 352301
rect 72402 352141 72493 352259
rect 72611 352141 72702 352259
rect 72402 351760 72702 352141
rect 74202 351760 74502 353061
rect 76002 351760 76302 353981
rect 77802 351760 78102 354901
rect 86802 355639 87102 355650
rect 86802 355521 86893 355639
rect 87011 355521 87102 355639
rect 86802 355479 87102 355521
rect 86802 355361 86893 355479
rect 87011 355361 87102 355479
rect 85002 354719 85302 354730
rect 85002 354601 85093 354719
rect 85211 354601 85302 354719
rect 85002 354559 85302 354601
rect 85002 354441 85093 354559
rect 85211 354441 85302 354559
rect 83202 353799 83502 353810
rect 83202 353681 83293 353799
rect 83411 353681 83502 353799
rect 83202 353639 83502 353681
rect 83202 353521 83293 353639
rect 83411 353521 83502 353639
rect 81402 352879 81702 352890
rect 81402 352761 81493 352879
rect 81611 352761 81702 352879
rect 81402 352719 81702 352761
rect 81402 352601 81493 352719
rect 81611 352601 81702 352719
rect 81402 351760 81702 352601
rect 83202 351760 83502 353521
rect 85002 351760 85302 354441
rect 86802 351760 87102 355361
rect 95802 355179 96102 355650
rect 95802 355061 95893 355179
rect 96011 355061 96102 355179
rect 95802 355019 96102 355061
rect 95802 354901 95893 355019
rect 96011 354901 96102 355019
rect 94002 354259 94302 354730
rect 94002 354141 94093 354259
rect 94211 354141 94302 354259
rect 94002 354099 94302 354141
rect 94002 353981 94093 354099
rect 94211 353981 94302 354099
rect 92202 353339 92502 353810
rect 92202 353221 92293 353339
rect 92411 353221 92502 353339
rect 92202 353179 92502 353221
rect 92202 353061 92293 353179
rect 92411 353061 92502 353179
rect 90402 352419 90702 352890
rect 90402 352301 90493 352419
rect 90611 352301 90702 352419
rect 90402 352259 90702 352301
rect 90402 352141 90493 352259
rect 90611 352141 90702 352259
rect 90402 351760 90702 352141
rect 92202 351760 92502 353061
rect 94002 351760 94302 353981
rect 95802 351760 96102 354901
rect 104802 355639 105102 355650
rect 104802 355521 104893 355639
rect 105011 355521 105102 355639
rect 104802 355479 105102 355521
rect 104802 355361 104893 355479
rect 105011 355361 105102 355479
rect 103002 354719 103302 354730
rect 103002 354601 103093 354719
rect 103211 354601 103302 354719
rect 103002 354559 103302 354601
rect 103002 354441 103093 354559
rect 103211 354441 103302 354559
rect 101202 353799 101502 353810
rect 101202 353681 101293 353799
rect 101411 353681 101502 353799
rect 101202 353639 101502 353681
rect 101202 353521 101293 353639
rect 101411 353521 101502 353639
rect 99402 352879 99702 352890
rect 99402 352761 99493 352879
rect 99611 352761 99702 352879
rect 99402 352719 99702 352761
rect 99402 352601 99493 352719
rect 99611 352601 99702 352719
rect 99402 351760 99702 352601
rect 101202 351760 101502 353521
rect 103002 351760 103302 354441
rect 104802 351760 105102 355361
rect 113802 355179 114102 355650
rect 113802 355061 113893 355179
rect 114011 355061 114102 355179
rect 113802 355019 114102 355061
rect 113802 354901 113893 355019
rect 114011 354901 114102 355019
rect 112002 354259 112302 354730
rect 112002 354141 112093 354259
rect 112211 354141 112302 354259
rect 112002 354099 112302 354141
rect 112002 353981 112093 354099
rect 112211 353981 112302 354099
rect 110202 353339 110502 353810
rect 110202 353221 110293 353339
rect 110411 353221 110502 353339
rect 110202 353179 110502 353221
rect 110202 353061 110293 353179
rect 110411 353061 110502 353179
rect 108402 352419 108702 352890
rect 108402 352301 108493 352419
rect 108611 352301 108702 352419
rect 108402 352259 108702 352301
rect 108402 352141 108493 352259
rect 108611 352141 108702 352259
rect 108402 351760 108702 352141
rect 110202 351760 110502 353061
rect 112002 351760 112302 353981
rect 113802 351760 114102 354901
rect 122802 355639 123102 355650
rect 122802 355521 122893 355639
rect 123011 355521 123102 355639
rect 122802 355479 123102 355521
rect 122802 355361 122893 355479
rect 123011 355361 123102 355479
rect 121002 354719 121302 354730
rect 121002 354601 121093 354719
rect 121211 354601 121302 354719
rect 121002 354559 121302 354601
rect 121002 354441 121093 354559
rect 121211 354441 121302 354559
rect 119202 353799 119502 353810
rect 119202 353681 119293 353799
rect 119411 353681 119502 353799
rect 119202 353639 119502 353681
rect 119202 353521 119293 353639
rect 119411 353521 119502 353639
rect 117402 352879 117702 352890
rect 117402 352761 117493 352879
rect 117611 352761 117702 352879
rect 117402 352719 117702 352761
rect 117402 352601 117493 352719
rect 117611 352601 117702 352719
rect 117402 351760 117702 352601
rect 119202 351760 119502 353521
rect 121002 351760 121302 354441
rect 122802 351760 123102 355361
rect 131802 355179 132102 355650
rect 131802 355061 131893 355179
rect 132011 355061 132102 355179
rect 131802 355019 132102 355061
rect 131802 354901 131893 355019
rect 132011 354901 132102 355019
rect 130002 354259 130302 354730
rect 130002 354141 130093 354259
rect 130211 354141 130302 354259
rect 130002 354099 130302 354141
rect 130002 353981 130093 354099
rect 130211 353981 130302 354099
rect 128202 353339 128502 353810
rect 128202 353221 128293 353339
rect 128411 353221 128502 353339
rect 128202 353179 128502 353221
rect 128202 353061 128293 353179
rect 128411 353061 128502 353179
rect 126402 352419 126702 352890
rect 126402 352301 126493 352419
rect 126611 352301 126702 352419
rect 126402 352259 126702 352301
rect 126402 352141 126493 352259
rect 126611 352141 126702 352259
rect 126402 351760 126702 352141
rect 128202 351760 128502 353061
rect 130002 351760 130302 353981
rect 131802 351760 132102 354901
rect 140802 355639 141102 355650
rect 140802 355521 140893 355639
rect 141011 355521 141102 355639
rect 140802 355479 141102 355521
rect 140802 355361 140893 355479
rect 141011 355361 141102 355479
rect 139002 354719 139302 354730
rect 139002 354601 139093 354719
rect 139211 354601 139302 354719
rect 139002 354559 139302 354601
rect 139002 354441 139093 354559
rect 139211 354441 139302 354559
rect 137202 353799 137502 353810
rect 137202 353681 137293 353799
rect 137411 353681 137502 353799
rect 137202 353639 137502 353681
rect 137202 353521 137293 353639
rect 137411 353521 137502 353639
rect 135402 352879 135702 352890
rect 135402 352761 135493 352879
rect 135611 352761 135702 352879
rect 135402 352719 135702 352761
rect 135402 352601 135493 352719
rect 135611 352601 135702 352719
rect 135402 351760 135702 352601
rect 137202 351760 137502 353521
rect 139002 351760 139302 354441
rect 140802 351760 141102 355361
rect 149802 355179 150102 355650
rect 149802 355061 149893 355179
rect 150011 355061 150102 355179
rect 149802 355019 150102 355061
rect 149802 354901 149893 355019
rect 150011 354901 150102 355019
rect 148002 354259 148302 354730
rect 148002 354141 148093 354259
rect 148211 354141 148302 354259
rect 148002 354099 148302 354141
rect 148002 353981 148093 354099
rect 148211 353981 148302 354099
rect 146202 353339 146502 353810
rect 146202 353221 146293 353339
rect 146411 353221 146502 353339
rect 146202 353179 146502 353221
rect 146202 353061 146293 353179
rect 146411 353061 146502 353179
rect 144402 352419 144702 352890
rect 144402 352301 144493 352419
rect 144611 352301 144702 352419
rect 144402 352259 144702 352301
rect 144402 352141 144493 352259
rect 144611 352141 144702 352259
rect 144402 351760 144702 352141
rect 146202 351760 146502 353061
rect 148002 351760 148302 353981
rect 149802 351760 150102 354901
rect 158802 355639 159102 355650
rect 158802 355521 158893 355639
rect 159011 355521 159102 355639
rect 158802 355479 159102 355521
rect 158802 355361 158893 355479
rect 159011 355361 159102 355479
rect 157002 354719 157302 354730
rect 157002 354601 157093 354719
rect 157211 354601 157302 354719
rect 157002 354559 157302 354601
rect 157002 354441 157093 354559
rect 157211 354441 157302 354559
rect 155202 353799 155502 353810
rect 155202 353681 155293 353799
rect 155411 353681 155502 353799
rect 155202 353639 155502 353681
rect 155202 353521 155293 353639
rect 155411 353521 155502 353639
rect 153402 352879 153702 352890
rect 153402 352761 153493 352879
rect 153611 352761 153702 352879
rect 153402 352719 153702 352761
rect 153402 352601 153493 352719
rect 153611 352601 153702 352719
rect 153402 351760 153702 352601
rect 155202 351760 155502 353521
rect 157002 351760 157302 354441
rect 158802 351760 159102 355361
rect 167802 355179 168102 355650
rect 167802 355061 167893 355179
rect 168011 355061 168102 355179
rect 167802 355019 168102 355061
rect 167802 354901 167893 355019
rect 168011 354901 168102 355019
rect 166002 354259 166302 354730
rect 166002 354141 166093 354259
rect 166211 354141 166302 354259
rect 166002 354099 166302 354141
rect 166002 353981 166093 354099
rect 166211 353981 166302 354099
rect 164202 353339 164502 353810
rect 164202 353221 164293 353339
rect 164411 353221 164502 353339
rect 164202 353179 164502 353221
rect 164202 353061 164293 353179
rect 164411 353061 164502 353179
rect 162402 352419 162702 352890
rect 162402 352301 162493 352419
rect 162611 352301 162702 352419
rect 162402 352259 162702 352301
rect 162402 352141 162493 352259
rect 162611 352141 162702 352259
rect 162402 351760 162702 352141
rect 164202 351760 164502 353061
rect 166002 351760 166302 353981
rect 167802 351760 168102 354901
rect 176802 355639 177102 355650
rect 176802 355521 176893 355639
rect 177011 355521 177102 355639
rect 176802 355479 177102 355521
rect 176802 355361 176893 355479
rect 177011 355361 177102 355479
rect 175002 354719 175302 354730
rect 175002 354601 175093 354719
rect 175211 354601 175302 354719
rect 175002 354559 175302 354601
rect 175002 354441 175093 354559
rect 175211 354441 175302 354559
rect 173202 353799 173502 353810
rect 173202 353681 173293 353799
rect 173411 353681 173502 353799
rect 173202 353639 173502 353681
rect 173202 353521 173293 353639
rect 173411 353521 173502 353639
rect 171402 352879 171702 352890
rect 171402 352761 171493 352879
rect 171611 352761 171702 352879
rect 171402 352719 171702 352761
rect 171402 352601 171493 352719
rect 171611 352601 171702 352719
rect 171402 351760 171702 352601
rect 173202 351760 173502 353521
rect 175002 351760 175302 354441
rect 176802 351760 177102 355361
rect 185802 355179 186102 355650
rect 185802 355061 185893 355179
rect 186011 355061 186102 355179
rect 185802 355019 186102 355061
rect 185802 354901 185893 355019
rect 186011 354901 186102 355019
rect 184002 354259 184302 354730
rect 184002 354141 184093 354259
rect 184211 354141 184302 354259
rect 184002 354099 184302 354141
rect 184002 353981 184093 354099
rect 184211 353981 184302 354099
rect 182202 353339 182502 353810
rect 182202 353221 182293 353339
rect 182411 353221 182502 353339
rect 182202 353179 182502 353221
rect 182202 353061 182293 353179
rect 182411 353061 182502 353179
rect 180402 352419 180702 352890
rect 180402 352301 180493 352419
rect 180611 352301 180702 352419
rect 180402 352259 180702 352301
rect 180402 352141 180493 352259
rect 180611 352141 180702 352259
rect 180402 351760 180702 352141
rect 182202 351760 182502 353061
rect 184002 351760 184302 353981
rect 185802 351760 186102 354901
rect 194802 355639 195102 355650
rect 194802 355521 194893 355639
rect 195011 355521 195102 355639
rect 194802 355479 195102 355521
rect 194802 355361 194893 355479
rect 195011 355361 195102 355479
rect 193002 354719 193302 354730
rect 193002 354601 193093 354719
rect 193211 354601 193302 354719
rect 193002 354559 193302 354601
rect 193002 354441 193093 354559
rect 193211 354441 193302 354559
rect 191202 353799 191502 353810
rect 191202 353681 191293 353799
rect 191411 353681 191502 353799
rect 191202 353639 191502 353681
rect 191202 353521 191293 353639
rect 191411 353521 191502 353639
rect 189402 352879 189702 352890
rect 189402 352761 189493 352879
rect 189611 352761 189702 352879
rect 189402 352719 189702 352761
rect 189402 352601 189493 352719
rect 189611 352601 189702 352719
rect 189402 351760 189702 352601
rect 191202 351760 191502 353521
rect 193002 351760 193302 354441
rect 194802 351760 195102 355361
rect 203802 355179 204102 355650
rect 203802 355061 203893 355179
rect 204011 355061 204102 355179
rect 203802 355019 204102 355061
rect 203802 354901 203893 355019
rect 204011 354901 204102 355019
rect 202002 354259 202302 354730
rect 202002 354141 202093 354259
rect 202211 354141 202302 354259
rect 202002 354099 202302 354141
rect 202002 353981 202093 354099
rect 202211 353981 202302 354099
rect 200202 353339 200502 353810
rect 200202 353221 200293 353339
rect 200411 353221 200502 353339
rect 200202 353179 200502 353221
rect 200202 353061 200293 353179
rect 200411 353061 200502 353179
rect 198402 352419 198702 352890
rect 198402 352301 198493 352419
rect 198611 352301 198702 352419
rect 198402 352259 198702 352301
rect 198402 352141 198493 352259
rect 198611 352141 198702 352259
rect 198402 351760 198702 352141
rect 200202 351760 200502 353061
rect 202002 351760 202302 353981
rect 203802 351760 204102 354901
rect 212802 355639 213102 355650
rect 212802 355521 212893 355639
rect 213011 355521 213102 355639
rect 212802 355479 213102 355521
rect 212802 355361 212893 355479
rect 213011 355361 213102 355479
rect 211002 354719 211302 354730
rect 211002 354601 211093 354719
rect 211211 354601 211302 354719
rect 211002 354559 211302 354601
rect 211002 354441 211093 354559
rect 211211 354441 211302 354559
rect 209202 353799 209502 353810
rect 209202 353681 209293 353799
rect 209411 353681 209502 353799
rect 209202 353639 209502 353681
rect 209202 353521 209293 353639
rect 209411 353521 209502 353639
rect 207402 352879 207702 352890
rect 207402 352761 207493 352879
rect 207611 352761 207702 352879
rect 207402 352719 207702 352761
rect 207402 352601 207493 352719
rect 207611 352601 207702 352719
rect 207402 351760 207702 352601
rect 209202 351760 209502 353521
rect 211002 351760 211302 354441
rect 212802 351760 213102 355361
rect 221802 355179 222102 355650
rect 221802 355061 221893 355179
rect 222011 355061 222102 355179
rect 221802 355019 222102 355061
rect 221802 354901 221893 355019
rect 222011 354901 222102 355019
rect 220002 354259 220302 354730
rect 220002 354141 220093 354259
rect 220211 354141 220302 354259
rect 220002 354099 220302 354141
rect 220002 353981 220093 354099
rect 220211 353981 220302 354099
rect 218202 353339 218502 353810
rect 218202 353221 218293 353339
rect 218411 353221 218502 353339
rect 218202 353179 218502 353221
rect 218202 353061 218293 353179
rect 218411 353061 218502 353179
rect 216402 352419 216702 352890
rect 216402 352301 216493 352419
rect 216611 352301 216702 352419
rect 216402 352259 216702 352301
rect 216402 352141 216493 352259
rect 216611 352141 216702 352259
rect 216402 351760 216702 352141
rect 218202 351760 218502 353061
rect 220002 351760 220302 353981
rect 221802 351760 222102 354901
rect 230802 355639 231102 355650
rect 230802 355521 230893 355639
rect 231011 355521 231102 355639
rect 230802 355479 231102 355521
rect 230802 355361 230893 355479
rect 231011 355361 231102 355479
rect 229002 354719 229302 354730
rect 229002 354601 229093 354719
rect 229211 354601 229302 354719
rect 229002 354559 229302 354601
rect 229002 354441 229093 354559
rect 229211 354441 229302 354559
rect 227202 353799 227502 353810
rect 227202 353681 227293 353799
rect 227411 353681 227502 353799
rect 227202 353639 227502 353681
rect 227202 353521 227293 353639
rect 227411 353521 227502 353639
rect 225402 352879 225702 352890
rect 225402 352761 225493 352879
rect 225611 352761 225702 352879
rect 225402 352719 225702 352761
rect 225402 352601 225493 352719
rect 225611 352601 225702 352719
rect 225402 351760 225702 352601
rect 227202 351760 227502 353521
rect 229002 351760 229302 354441
rect 230802 351760 231102 355361
rect 239802 355179 240102 355650
rect 239802 355061 239893 355179
rect 240011 355061 240102 355179
rect 239802 355019 240102 355061
rect 239802 354901 239893 355019
rect 240011 354901 240102 355019
rect 238002 354259 238302 354730
rect 238002 354141 238093 354259
rect 238211 354141 238302 354259
rect 238002 354099 238302 354141
rect 238002 353981 238093 354099
rect 238211 353981 238302 354099
rect 236202 353339 236502 353810
rect 236202 353221 236293 353339
rect 236411 353221 236502 353339
rect 236202 353179 236502 353221
rect 236202 353061 236293 353179
rect 236411 353061 236502 353179
rect 234402 352419 234702 352890
rect 234402 352301 234493 352419
rect 234611 352301 234702 352419
rect 234402 352259 234702 352301
rect 234402 352141 234493 352259
rect 234611 352141 234702 352259
rect 234402 351760 234702 352141
rect 236202 351760 236502 353061
rect 238002 351760 238302 353981
rect 239802 351760 240102 354901
rect 248802 355639 249102 355650
rect 248802 355521 248893 355639
rect 249011 355521 249102 355639
rect 248802 355479 249102 355521
rect 248802 355361 248893 355479
rect 249011 355361 249102 355479
rect 247002 354719 247302 354730
rect 247002 354601 247093 354719
rect 247211 354601 247302 354719
rect 247002 354559 247302 354601
rect 247002 354441 247093 354559
rect 247211 354441 247302 354559
rect 245202 353799 245502 353810
rect 245202 353681 245293 353799
rect 245411 353681 245502 353799
rect 245202 353639 245502 353681
rect 245202 353521 245293 353639
rect 245411 353521 245502 353639
rect 243402 352879 243702 352890
rect 243402 352761 243493 352879
rect 243611 352761 243702 352879
rect 243402 352719 243702 352761
rect 243402 352601 243493 352719
rect 243611 352601 243702 352719
rect 243402 351760 243702 352601
rect 245202 351760 245502 353521
rect 247002 351760 247302 354441
rect 248802 351760 249102 355361
rect 257802 355179 258102 355650
rect 257802 355061 257893 355179
rect 258011 355061 258102 355179
rect 257802 355019 258102 355061
rect 257802 354901 257893 355019
rect 258011 354901 258102 355019
rect 256002 354259 256302 354730
rect 256002 354141 256093 354259
rect 256211 354141 256302 354259
rect 256002 354099 256302 354141
rect 256002 353981 256093 354099
rect 256211 353981 256302 354099
rect 254202 353339 254502 353810
rect 254202 353221 254293 353339
rect 254411 353221 254502 353339
rect 254202 353179 254502 353221
rect 254202 353061 254293 353179
rect 254411 353061 254502 353179
rect 252402 352419 252702 352890
rect 252402 352301 252493 352419
rect 252611 352301 252702 352419
rect 252402 352259 252702 352301
rect 252402 352141 252493 352259
rect 252611 352141 252702 352259
rect 252402 351760 252702 352141
rect 254202 351760 254502 353061
rect 256002 351760 256302 353981
rect 257802 351760 258102 354901
rect 266802 355639 267102 355650
rect 266802 355521 266893 355639
rect 267011 355521 267102 355639
rect 266802 355479 267102 355521
rect 266802 355361 266893 355479
rect 267011 355361 267102 355479
rect 265002 354719 265302 354730
rect 265002 354601 265093 354719
rect 265211 354601 265302 354719
rect 265002 354559 265302 354601
rect 265002 354441 265093 354559
rect 265211 354441 265302 354559
rect 263202 353799 263502 353810
rect 263202 353681 263293 353799
rect 263411 353681 263502 353799
rect 263202 353639 263502 353681
rect 263202 353521 263293 353639
rect 263411 353521 263502 353639
rect 261402 352879 261702 352890
rect 261402 352761 261493 352879
rect 261611 352761 261702 352879
rect 261402 352719 261702 352761
rect 261402 352601 261493 352719
rect 261611 352601 261702 352719
rect 261402 351760 261702 352601
rect 263202 351760 263502 353521
rect 265002 351760 265302 354441
rect 266802 351760 267102 355361
rect 275802 355179 276102 355650
rect 275802 355061 275893 355179
rect 276011 355061 276102 355179
rect 275802 355019 276102 355061
rect 275802 354901 275893 355019
rect 276011 354901 276102 355019
rect 274002 354259 274302 354730
rect 274002 354141 274093 354259
rect 274211 354141 274302 354259
rect 274002 354099 274302 354141
rect 274002 353981 274093 354099
rect 274211 353981 274302 354099
rect 272202 353339 272502 353810
rect 272202 353221 272293 353339
rect 272411 353221 272502 353339
rect 272202 353179 272502 353221
rect 272202 353061 272293 353179
rect 272411 353061 272502 353179
rect 270402 352419 270702 352890
rect 270402 352301 270493 352419
rect 270611 352301 270702 352419
rect 270402 352259 270702 352301
rect 270402 352141 270493 352259
rect 270611 352141 270702 352259
rect 270402 351760 270702 352141
rect 272202 351760 272502 353061
rect 274002 351760 274302 353981
rect 275802 351760 276102 354901
rect 284802 355639 285102 355650
rect 284802 355521 284893 355639
rect 285011 355521 285102 355639
rect 284802 355479 285102 355521
rect 284802 355361 284893 355479
rect 285011 355361 285102 355479
rect 283002 354719 283302 354730
rect 283002 354601 283093 354719
rect 283211 354601 283302 354719
rect 283002 354559 283302 354601
rect 283002 354441 283093 354559
rect 283211 354441 283302 354559
rect 281202 353799 281502 353810
rect 281202 353681 281293 353799
rect 281411 353681 281502 353799
rect 281202 353639 281502 353681
rect 281202 353521 281293 353639
rect 281411 353521 281502 353639
rect 279402 352879 279702 352890
rect 279402 352761 279493 352879
rect 279611 352761 279702 352879
rect 279402 352719 279702 352761
rect 279402 352601 279493 352719
rect 279611 352601 279702 352719
rect 279402 351760 279702 352601
rect 281202 351760 281502 353521
rect 283002 351760 283302 354441
rect 284802 351760 285102 355361
rect 295880 355639 296180 355650
rect 295880 355521 295971 355639
rect 296089 355521 296180 355639
rect 295880 355479 296180 355521
rect 295880 355361 295971 355479
rect 296089 355361 296180 355479
rect 295420 355179 295720 355190
rect 295420 355061 295511 355179
rect 295629 355061 295720 355179
rect 295420 355019 295720 355061
rect 295420 354901 295511 355019
rect 295629 354901 295720 355019
rect 294960 354719 295260 354730
rect 294960 354601 295051 354719
rect 295169 354601 295260 354719
rect 294960 354559 295260 354601
rect 294960 354441 295051 354559
rect 295169 354441 295260 354559
rect 294500 354259 294800 354270
rect 294500 354141 294591 354259
rect 294709 354141 294800 354259
rect 294500 354099 294800 354141
rect 294500 353981 294591 354099
rect 294709 353981 294800 354099
rect 290202 353339 290502 353810
rect 294040 353799 294340 353810
rect 294040 353681 294131 353799
rect 294249 353681 294340 353799
rect 294040 353639 294340 353681
rect 294040 353521 294131 353639
rect 294249 353521 294340 353639
rect 290202 353221 290293 353339
rect 290411 353221 290502 353339
rect 290202 353179 290502 353221
rect 290202 353061 290293 353179
rect 290411 353061 290502 353179
rect 288402 352419 288702 352890
rect 288402 352301 288493 352419
rect 288611 352301 288702 352419
rect 288402 352259 288702 352301
rect 288402 352141 288493 352259
rect 288611 352141 288702 352259
rect 288402 351760 288702 352141
rect 290202 351760 290502 353061
rect 293580 353339 293880 353350
rect 293580 353221 293671 353339
rect 293789 353221 293880 353339
rect 293580 353179 293880 353221
rect 293580 353061 293671 353179
rect 293789 353061 293880 353179
rect 293120 352879 293420 352890
rect 293120 352761 293211 352879
rect 293329 352761 293420 352879
rect 293120 352719 293420 352761
rect 293120 352601 293211 352719
rect 293329 352601 293420 352719
rect 292660 352419 292960 352430
rect 292660 352301 292751 352419
rect 292869 352301 292960 352419
rect 292660 352259 292960 352301
rect 292660 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 343109 -907 343227
rect -789 343109 -698 343227
rect -998 343067 -698 343109
rect -998 342949 -907 343067
rect -789 342949 -698 343067
rect -998 325227 -698 342949
rect -998 325109 -907 325227
rect -789 325109 -698 325227
rect -998 325067 -698 325109
rect -998 324949 -907 325067
rect -789 324949 -698 325067
rect -998 307227 -698 324949
rect -998 307109 -907 307227
rect -789 307109 -698 307227
rect -998 307067 -698 307109
rect -998 306949 -907 307067
rect -789 306949 -698 307067
rect -998 289227 -698 306949
rect -998 289109 -907 289227
rect -789 289109 -698 289227
rect -998 289067 -698 289109
rect -998 288949 -907 289067
rect -789 288949 -698 289067
rect -998 271227 -698 288949
rect -998 271109 -907 271227
rect -789 271109 -698 271227
rect -998 271067 -698 271109
rect -998 270949 -907 271067
rect -789 270949 -698 271067
rect -998 253227 -698 270949
rect -998 253109 -907 253227
rect -789 253109 -698 253227
rect -998 253067 -698 253109
rect -998 252949 -907 253067
rect -789 252949 -698 253067
rect -998 235227 -698 252949
rect -998 235109 -907 235227
rect -789 235109 -698 235227
rect -998 235067 -698 235109
rect -998 234949 -907 235067
rect -789 234949 -698 235067
rect -998 217227 -698 234949
rect -998 217109 -907 217227
rect -789 217109 -698 217227
rect -998 217067 -698 217109
rect -998 216949 -907 217067
rect -789 216949 -698 217067
rect -998 199227 -698 216949
rect -998 199109 -907 199227
rect -789 199109 -698 199227
rect -998 199067 -698 199109
rect -998 198949 -907 199067
rect -789 198949 -698 199067
rect -998 181227 -698 198949
rect -998 181109 -907 181227
rect -789 181109 -698 181227
rect -998 181067 -698 181109
rect -998 180949 -907 181067
rect -789 180949 -698 181067
rect -998 163227 -698 180949
rect -998 163109 -907 163227
rect -789 163109 -698 163227
rect -998 163067 -698 163109
rect -998 162949 -907 163067
rect -789 162949 -698 163067
rect -998 145227 -698 162949
rect -998 145109 -907 145227
rect -789 145109 -698 145227
rect -998 145067 -698 145109
rect -998 144949 -907 145067
rect -789 144949 -698 145067
rect -998 127227 -698 144949
rect -998 127109 -907 127227
rect -789 127109 -698 127227
rect -998 127067 -698 127109
rect -998 126949 -907 127067
rect -789 126949 -698 127067
rect -998 109227 -698 126949
rect -998 109109 -907 109227
rect -789 109109 -698 109227
rect -998 109067 -698 109109
rect -998 108949 -907 109067
rect -789 108949 -698 109067
rect -998 91227 -698 108949
rect -998 91109 -907 91227
rect -789 91109 -698 91227
rect -998 91067 -698 91109
rect -998 90949 -907 91067
rect -789 90949 -698 91067
rect -998 73227 -698 90949
rect -998 73109 -907 73227
rect -789 73109 -698 73227
rect -998 73067 -698 73109
rect -998 72949 -907 73067
rect -789 72949 -698 73067
rect -998 55227 -698 72949
rect -998 55109 -907 55227
rect -789 55109 -698 55227
rect -998 55067 -698 55109
rect -998 54949 -907 55067
rect -789 54949 -698 55067
rect -998 37227 -698 54949
rect -998 37109 -907 37227
rect -789 37109 -698 37227
rect -998 37067 -698 37109
rect -998 36949 -907 37067
rect -789 36949 -698 37067
rect -998 19227 -698 36949
rect -998 19109 -907 19227
rect -789 19109 -698 19227
rect -998 19067 -698 19109
rect -998 18949 -907 19067
rect -789 18949 -698 19067
rect -998 1227 -698 18949
rect -998 1109 -907 1227
rect -789 1109 -698 1227
rect -998 1067 -698 1109
rect -998 949 -907 1067
rect -789 949 -698 1067
rect -998 -173 -698 949
rect 292660 343227 292960 352141
rect 292660 343109 292751 343227
rect 292869 343109 292960 343227
rect 292660 343067 292960 343109
rect 292660 342949 292751 343067
rect 292869 342949 292960 343067
rect 292660 325227 292960 342949
rect 292660 325109 292751 325227
rect 292869 325109 292960 325227
rect 292660 325067 292960 325109
rect 292660 324949 292751 325067
rect 292869 324949 292960 325067
rect 292660 307227 292960 324949
rect 292660 307109 292751 307227
rect 292869 307109 292960 307227
rect 292660 307067 292960 307109
rect 292660 306949 292751 307067
rect 292869 306949 292960 307067
rect 292660 289227 292960 306949
rect 292660 289109 292751 289227
rect 292869 289109 292960 289227
rect 292660 289067 292960 289109
rect 292660 288949 292751 289067
rect 292869 288949 292960 289067
rect 292660 271227 292960 288949
rect 292660 271109 292751 271227
rect 292869 271109 292960 271227
rect 292660 271067 292960 271109
rect 292660 270949 292751 271067
rect 292869 270949 292960 271067
rect 292660 253227 292960 270949
rect 292660 253109 292751 253227
rect 292869 253109 292960 253227
rect 292660 253067 292960 253109
rect 292660 252949 292751 253067
rect 292869 252949 292960 253067
rect 292660 235227 292960 252949
rect 292660 235109 292751 235227
rect 292869 235109 292960 235227
rect 292660 235067 292960 235109
rect 292660 234949 292751 235067
rect 292869 234949 292960 235067
rect 292660 217227 292960 234949
rect 292660 217109 292751 217227
rect 292869 217109 292960 217227
rect 292660 217067 292960 217109
rect 292660 216949 292751 217067
rect 292869 216949 292960 217067
rect 292660 199227 292960 216949
rect 292660 199109 292751 199227
rect 292869 199109 292960 199227
rect 292660 199067 292960 199109
rect 292660 198949 292751 199067
rect 292869 198949 292960 199067
rect 292660 181227 292960 198949
rect 292660 181109 292751 181227
rect 292869 181109 292960 181227
rect 292660 181067 292960 181109
rect 292660 180949 292751 181067
rect 292869 180949 292960 181067
rect 292660 163227 292960 180949
rect 292660 163109 292751 163227
rect 292869 163109 292960 163227
rect 292660 163067 292960 163109
rect 292660 162949 292751 163067
rect 292869 162949 292960 163067
rect 292660 145227 292960 162949
rect 292660 145109 292751 145227
rect 292869 145109 292960 145227
rect 292660 145067 292960 145109
rect 292660 144949 292751 145067
rect 292869 144949 292960 145067
rect 292660 127227 292960 144949
rect 292660 127109 292751 127227
rect 292869 127109 292960 127227
rect 292660 127067 292960 127109
rect 292660 126949 292751 127067
rect 292869 126949 292960 127067
rect 292660 109227 292960 126949
rect 292660 109109 292751 109227
rect 292869 109109 292960 109227
rect 292660 109067 292960 109109
rect 292660 108949 292751 109067
rect 292869 108949 292960 109067
rect 292660 91227 292960 108949
rect 292660 91109 292751 91227
rect 292869 91109 292960 91227
rect 292660 91067 292960 91109
rect 292660 90949 292751 91067
rect 292869 90949 292960 91067
rect 292660 73227 292960 90949
rect 292660 73109 292751 73227
rect 292869 73109 292960 73227
rect 292660 73067 292960 73109
rect 292660 72949 292751 73067
rect 292869 72949 292960 73067
rect 292660 55227 292960 72949
rect 292660 55109 292751 55227
rect 292869 55109 292960 55227
rect 292660 55067 292960 55109
rect 292660 54949 292751 55067
rect 292869 54949 292960 55067
rect 292660 37227 292960 54949
rect 292660 37109 292751 37227
rect 292869 37109 292960 37227
rect 292660 37067 292960 37109
rect 292660 36949 292751 37067
rect 292869 36949 292960 37067
rect 292660 19227 292960 36949
rect 292660 19109 292751 19227
rect 292869 19109 292960 19227
rect 292660 19067 292960 19109
rect 292660 18949 292751 19067
rect 292869 18949 292960 19067
rect 292660 1227 292960 18949
rect 292660 1109 292751 1227
rect 292869 1109 292960 1227
rect 292660 1067 292960 1109
rect 292660 949 292751 1067
rect 292869 949 292960 1067
rect -998 -291 -907 -173
rect -789 -291 -698 -173
rect -998 -333 -698 -291
rect -998 -451 -907 -333
rect -789 -451 -698 -333
rect -998 -462 -698 -451
rect 402 -173 702 240
rect 402 -291 493 -173
rect 611 -291 702 -173
rect 402 -333 702 -291
rect 402 -451 493 -333
rect 611 -451 702 -333
rect -1458 -751 -1367 -633
rect -1249 -751 -1158 -633
rect -1458 -793 -1158 -751
rect -1458 -911 -1367 -793
rect -1249 -911 -1158 -793
rect -1458 -922 -1158 -911
rect 402 -922 702 -451
rect -1918 -1211 -1827 -1093
rect -1709 -1211 -1618 -1093
rect -1918 -1253 -1618 -1211
rect -1918 -1371 -1827 -1253
rect -1709 -1371 -1618 -1253
rect -1918 -1382 -1618 -1371
rect 2202 -1093 2502 240
rect 2202 -1211 2293 -1093
rect 2411 -1211 2502 -1093
rect 2202 -1253 2502 -1211
rect 2202 -1371 2293 -1253
rect 2411 -1371 2502 -1253
rect -2378 -1671 -2287 -1553
rect -2169 -1671 -2078 -1553
rect -2378 -1713 -2078 -1671
rect -2378 -1831 -2287 -1713
rect -2169 -1831 -2078 -1713
rect -2378 -1842 -2078 -1831
rect 2202 -1842 2502 -1371
rect -2838 -2131 -2747 -2013
rect -2629 -2131 -2538 -2013
rect -2838 -2173 -2538 -2131
rect -2838 -2291 -2747 -2173
rect -2629 -2291 -2538 -2173
rect -2838 -2302 -2538 -2291
rect 4002 -2013 4302 240
rect 4002 -2131 4093 -2013
rect 4211 -2131 4302 -2013
rect 4002 -2173 4302 -2131
rect 4002 -2291 4093 -2173
rect 4211 -2291 4302 -2173
rect -3298 -2591 -3207 -2473
rect -3089 -2591 -2998 -2473
rect -3298 -2633 -2998 -2591
rect -3298 -2751 -3207 -2633
rect -3089 -2751 -2998 -2633
rect -3298 -2762 -2998 -2751
rect 4002 -2762 4302 -2291
rect -3758 -3051 -3667 -2933
rect -3549 -3051 -3458 -2933
rect -3758 -3093 -3458 -3051
rect -3758 -3211 -3667 -3093
rect -3549 -3211 -3458 -3093
rect -3758 -3222 -3458 -3211
rect 5802 -2933 6102 240
rect 9402 -633 9702 240
rect 9402 -751 9493 -633
rect 9611 -751 9702 -633
rect 9402 -793 9702 -751
rect 9402 -911 9493 -793
rect 9611 -911 9702 -793
rect 9402 -922 9702 -911
rect 11202 -1553 11502 240
rect 11202 -1671 11293 -1553
rect 11411 -1671 11502 -1553
rect 11202 -1713 11502 -1671
rect 11202 -1831 11293 -1713
rect 11411 -1831 11502 -1713
rect 11202 -1842 11502 -1831
rect 13002 -2473 13302 240
rect 13002 -2591 13093 -2473
rect 13211 -2591 13302 -2473
rect 13002 -2633 13302 -2591
rect 13002 -2751 13093 -2633
rect 13211 -2751 13302 -2633
rect 13002 -2762 13302 -2751
rect 5802 -3051 5893 -2933
rect 6011 -3051 6102 -2933
rect 5802 -3093 6102 -3051
rect 5802 -3211 5893 -3093
rect 6011 -3211 6102 -3093
rect -4218 -3511 -4127 -3393
rect -4009 -3511 -3918 -3393
rect -4218 -3553 -3918 -3511
rect -4218 -3671 -4127 -3553
rect -4009 -3671 -3918 -3553
rect -4218 -3682 -3918 -3671
rect 5802 -3682 6102 -3211
rect 14802 -3393 15102 240
rect 18402 -173 18702 240
rect 18402 -291 18493 -173
rect 18611 -291 18702 -173
rect 18402 -333 18702 -291
rect 18402 -451 18493 -333
rect 18611 -451 18702 -333
rect 18402 -922 18702 -451
rect 20202 -1093 20502 240
rect 20202 -1211 20293 -1093
rect 20411 -1211 20502 -1093
rect 20202 -1253 20502 -1211
rect 20202 -1371 20293 -1253
rect 20411 -1371 20502 -1253
rect 20202 -1842 20502 -1371
rect 22002 -2013 22302 240
rect 22002 -2131 22093 -2013
rect 22211 -2131 22302 -2013
rect 22002 -2173 22302 -2131
rect 22002 -2291 22093 -2173
rect 22211 -2291 22302 -2173
rect 22002 -2762 22302 -2291
rect 14802 -3511 14893 -3393
rect 15011 -3511 15102 -3393
rect 14802 -3553 15102 -3511
rect 14802 -3671 14893 -3553
rect 15011 -3671 15102 -3553
rect 14802 -3682 15102 -3671
rect 23802 -2933 24102 240
rect 27402 -633 27702 240
rect 27402 -751 27493 -633
rect 27611 -751 27702 -633
rect 27402 -793 27702 -751
rect 27402 -911 27493 -793
rect 27611 -911 27702 -793
rect 27402 -922 27702 -911
rect 29202 -1553 29502 240
rect 29202 -1671 29293 -1553
rect 29411 -1671 29502 -1553
rect 29202 -1713 29502 -1671
rect 29202 -1831 29293 -1713
rect 29411 -1831 29502 -1713
rect 29202 -1842 29502 -1831
rect 31002 -2473 31302 240
rect 31002 -2591 31093 -2473
rect 31211 -2591 31302 -2473
rect 31002 -2633 31302 -2591
rect 31002 -2751 31093 -2633
rect 31211 -2751 31302 -2633
rect 31002 -2762 31302 -2751
rect 23802 -3051 23893 -2933
rect 24011 -3051 24102 -2933
rect 23802 -3093 24102 -3051
rect 23802 -3211 23893 -3093
rect 24011 -3211 24102 -3093
rect 23802 -3682 24102 -3211
rect 32802 -3393 33102 240
rect 36402 -173 36702 240
rect 36402 -291 36493 -173
rect 36611 -291 36702 -173
rect 36402 -333 36702 -291
rect 36402 -451 36493 -333
rect 36611 -451 36702 -333
rect 36402 -922 36702 -451
rect 38202 -1093 38502 240
rect 38202 -1211 38293 -1093
rect 38411 -1211 38502 -1093
rect 38202 -1253 38502 -1211
rect 38202 -1371 38293 -1253
rect 38411 -1371 38502 -1253
rect 38202 -1842 38502 -1371
rect 40002 -2013 40302 240
rect 40002 -2131 40093 -2013
rect 40211 -2131 40302 -2013
rect 40002 -2173 40302 -2131
rect 40002 -2291 40093 -2173
rect 40211 -2291 40302 -2173
rect 40002 -2762 40302 -2291
rect 32802 -3511 32893 -3393
rect 33011 -3511 33102 -3393
rect 32802 -3553 33102 -3511
rect 32802 -3671 32893 -3553
rect 33011 -3671 33102 -3553
rect 32802 -3682 33102 -3671
rect 41802 -2933 42102 240
rect 45402 -633 45702 240
rect 45402 -751 45493 -633
rect 45611 -751 45702 -633
rect 45402 -793 45702 -751
rect 45402 -911 45493 -793
rect 45611 -911 45702 -793
rect 45402 -922 45702 -911
rect 47202 -1553 47502 240
rect 47202 -1671 47293 -1553
rect 47411 -1671 47502 -1553
rect 47202 -1713 47502 -1671
rect 47202 -1831 47293 -1713
rect 47411 -1831 47502 -1713
rect 47202 -1842 47502 -1831
rect 49002 -2473 49302 240
rect 49002 -2591 49093 -2473
rect 49211 -2591 49302 -2473
rect 49002 -2633 49302 -2591
rect 49002 -2751 49093 -2633
rect 49211 -2751 49302 -2633
rect 49002 -2762 49302 -2751
rect 41802 -3051 41893 -2933
rect 42011 -3051 42102 -2933
rect 41802 -3093 42102 -3051
rect 41802 -3211 41893 -3093
rect 42011 -3211 42102 -3093
rect 41802 -3682 42102 -3211
rect 50802 -3393 51102 240
rect 54402 -173 54702 240
rect 54402 -291 54493 -173
rect 54611 -291 54702 -173
rect 54402 -333 54702 -291
rect 54402 -451 54493 -333
rect 54611 -451 54702 -333
rect 54402 -922 54702 -451
rect 56202 -1093 56502 240
rect 56202 -1211 56293 -1093
rect 56411 -1211 56502 -1093
rect 56202 -1253 56502 -1211
rect 56202 -1371 56293 -1253
rect 56411 -1371 56502 -1253
rect 56202 -1842 56502 -1371
rect 58002 -2013 58302 240
rect 58002 -2131 58093 -2013
rect 58211 -2131 58302 -2013
rect 58002 -2173 58302 -2131
rect 58002 -2291 58093 -2173
rect 58211 -2291 58302 -2173
rect 58002 -2762 58302 -2291
rect 50802 -3511 50893 -3393
rect 51011 -3511 51102 -3393
rect 50802 -3553 51102 -3511
rect 50802 -3671 50893 -3553
rect 51011 -3671 51102 -3553
rect 50802 -3682 51102 -3671
rect 59802 -2933 60102 240
rect 63402 -633 63702 240
rect 63402 -751 63493 -633
rect 63611 -751 63702 -633
rect 63402 -793 63702 -751
rect 63402 -911 63493 -793
rect 63611 -911 63702 -793
rect 63402 -922 63702 -911
rect 65202 -1553 65502 240
rect 65202 -1671 65293 -1553
rect 65411 -1671 65502 -1553
rect 65202 -1713 65502 -1671
rect 65202 -1831 65293 -1713
rect 65411 -1831 65502 -1713
rect 65202 -1842 65502 -1831
rect 67002 -2473 67302 240
rect 67002 -2591 67093 -2473
rect 67211 -2591 67302 -2473
rect 67002 -2633 67302 -2591
rect 67002 -2751 67093 -2633
rect 67211 -2751 67302 -2633
rect 67002 -2762 67302 -2751
rect 59802 -3051 59893 -2933
rect 60011 -3051 60102 -2933
rect 59802 -3093 60102 -3051
rect 59802 -3211 59893 -3093
rect 60011 -3211 60102 -3093
rect 59802 -3682 60102 -3211
rect 68802 -3393 69102 240
rect 72402 -173 72702 240
rect 72402 -291 72493 -173
rect 72611 -291 72702 -173
rect 72402 -333 72702 -291
rect 72402 -451 72493 -333
rect 72611 -451 72702 -333
rect 72402 -922 72702 -451
rect 74202 -1093 74502 240
rect 74202 -1211 74293 -1093
rect 74411 -1211 74502 -1093
rect 74202 -1253 74502 -1211
rect 74202 -1371 74293 -1253
rect 74411 -1371 74502 -1253
rect 74202 -1842 74502 -1371
rect 76002 -2013 76302 240
rect 76002 -2131 76093 -2013
rect 76211 -2131 76302 -2013
rect 76002 -2173 76302 -2131
rect 76002 -2291 76093 -2173
rect 76211 -2291 76302 -2173
rect 76002 -2762 76302 -2291
rect 68802 -3511 68893 -3393
rect 69011 -3511 69102 -3393
rect 68802 -3553 69102 -3511
rect 68802 -3671 68893 -3553
rect 69011 -3671 69102 -3553
rect 68802 -3682 69102 -3671
rect 77802 -2933 78102 240
rect 81402 -633 81702 240
rect 81402 -751 81493 -633
rect 81611 -751 81702 -633
rect 81402 -793 81702 -751
rect 81402 -911 81493 -793
rect 81611 -911 81702 -793
rect 81402 -922 81702 -911
rect 83202 -1553 83502 240
rect 83202 -1671 83293 -1553
rect 83411 -1671 83502 -1553
rect 83202 -1713 83502 -1671
rect 83202 -1831 83293 -1713
rect 83411 -1831 83502 -1713
rect 83202 -1842 83502 -1831
rect 85002 -2473 85302 240
rect 85002 -2591 85093 -2473
rect 85211 -2591 85302 -2473
rect 85002 -2633 85302 -2591
rect 85002 -2751 85093 -2633
rect 85211 -2751 85302 -2633
rect 85002 -2762 85302 -2751
rect 77802 -3051 77893 -2933
rect 78011 -3051 78102 -2933
rect 77802 -3093 78102 -3051
rect 77802 -3211 77893 -3093
rect 78011 -3211 78102 -3093
rect 77802 -3682 78102 -3211
rect 86802 -3393 87102 240
rect 90402 -173 90702 240
rect 90402 -291 90493 -173
rect 90611 -291 90702 -173
rect 90402 -333 90702 -291
rect 90402 -451 90493 -333
rect 90611 -451 90702 -333
rect 90402 -922 90702 -451
rect 92202 -1093 92502 240
rect 92202 -1211 92293 -1093
rect 92411 -1211 92502 -1093
rect 92202 -1253 92502 -1211
rect 92202 -1371 92293 -1253
rect 92411 -1371 92502 -1253
rect 92202 -1842 92502 -1371
rect 94002 -2013 94302 240
rect 94002 -2131 94093 -2013
rect 94211 -2131 94302 -2013
rect 94002 -2173 94302 -2131
rect 94002 -2291 94093 -2173
rect 94211 -2291 94302 -2173
rect 94002 -2762 94302 -2291
rect 86802 -3511 86893 -3393
rect 87011 -3511 87102 -3393
rect 86802 -3553 87102 -3511
rect 86802 -3671 86893 -3553
rect 87011 -3671 87102 -3553
rect 86802 -3682 87102 -3671
rect 95802 -2933 96102 240
rect 99402 -633 99702 240
rect 99402 -751 99493 -633
rect 99611 -751 99702 -633
rect 99402 -793 99702 -751
rect 99402 -911 99493 -793
rect 99611 -911 99702 -793
rect 99402 -922 99702 -911
rect 101202 -1553 101502 240
rect 101202 -1671 101293 -1553
rect 101411 -1671 101502 -1553
rect 101202 -1713 101502 -1671
rect 101202 -1831 101293 -1713
rect 101411 -1831 101502 -1713
rect 101202 -1842 101502 -1831
rect 103002 -2473 103302 240
rect 103002 -2591 103093 -2473
rect 103211 -2591 103302 -2473
rect 103002 -2633 103302 -2591
rect 103002 -2751 103093 -2633
rect 103211 -2751 103302 -2633
rect 103002 -2762 103302 -2751
rect 95802 -3051 95893 -2933
rect 96011 -3051 96102 -2933
rect 95802 -3093 96102 -3051
rect 95802 -3211 95893 -3093
rect 96011 -3211 96102 -3093
rect 95802 -3682 96102 -3211
rect 104802 -3393 105102 240
rect 108402 -173 108702 240
rect 108402 -291 108493 -173
rect 108611 -291 108702 -173
rect 108402 -333 108702 -291
rect 108402 -451 108493 -333
rect 108611 -451 108702 -333
rect 108402 -922 108702 -451
rect 110202 -1093 110502 240
rect 110202 -1211 110293 -1093
rect 110411 -1211 110502 -1093
rect 110202 -1253 110502 -1211
rect 110202 -1371 110293 -1253
rect 110411 -1371 110502 -1253
rect 110202 -1842 110502 -1371
rect 112002 -2013 112302 240
rect 112002 -2131 112093 -2013
rect 112211 -2131 112302 -2013
rect 112002 -2173 112302 -2131
rect 112002 -2291 112093 -2173
rect 112211 -2291 112302 -2173
rect 112002 -2762 112302 -2291
rect 104802 -3511 104893 -3393
rect 105011 -3511 105102 -3393
rect 104802 -3553 105102 -3511
rect 104802 -3671 104893 -3553
rect 105011 -3671 105102 -3553
rect 104802 -3682 105102 -3671
rect 113802 -2933 114102 240
rect 117402 -633 117702 240
rect 117402 -751 117493 -633
rect 117611 -751 117702 -633
rect 117402 -793 117702 -751
rect 117402 -911 117493 -793
rect 117611 -911 117702 -793
rect 117402 -922 117702 -911
rect 119202 -1553 119502 240
rect 119202 -1671 119293 -1553
rect 119411 -1671 119502 -1553
rect 119202 -1713 119502 -1671
rect 119202 -1831 119293 -1713
rect 119411 -1831 119502 -1713
rect 119202 -1842 119502 -1831
rect 121002 -2473 121302 240
rect 121002 -2591 121093 -2473
rect 121211 -2591 121302 -2473
rect 121002 -2633 121302 -2591
rect 121002 -2751 121093 -2633
rect 121211 -2751 121302 -2633
rect 121002 -2762 121302 -2751
rect 113802 -3051 113893 -2933
rect 114011 -3051 114102 -2933
rect 113802 -3093 114102 -3051
rect 113802 -3211 113893 -3093
rect 114011 -3211 114102 -3093
rect 113802 -3682 114102 -3211
rect 122802 -3393 123102 240
rect 126402 -173 126702 240
rect 126402 -291 126493 -173
rect 126611 -291 126702 -173
rect 126402 -333 126702 -291
rect 126402 -451 126493 -333
rect 126611 -451 126702 -333
rect 126402 -922 126702 -451
rect 128202 -1093 128502 240
rect 128202 -1211 128293 -1093
rect 128411 -1211 128502 -1093
rect 128202 -1253 128502 -1211
rect 128202 -1371 128293 -1253
rect 128411 -1371 128502 -1253
rect 128202 -1842 128502 -1371
rect 130002 -2013 130302 240
rect 130002 -2131 130093 -2013
rect 130211 -2131 130302 -2013
rect 130002 -2173 130302 -2131
rect 130002 -2291 130093 -2173
rect 130211 -2291 130302 -2173
rect 130002 -2762 130302 -2291
rect 122802 -3511 122893 -3393
rect 123011 -3511 123102 -3393
rect 122802 -3553 123102 -3511
rect 122802 -3671 122893 -3553
rect 123011 -3671 123102 -3553
rect 122802 -3682 123102 -3671
rect 131802 -2933 132102 240
rect 135402 -633 135702 240
rect 135402 -751 135493 -633
rect 135611 -751 135702 -633
rect 135402 -793 135702 -751
rect 135402 -911 135493 -793
rect 135611 -911 135702 -793
rect 135402 -922 135702 -911
rect 137202 -1553 137502 240
rect 137202 -1671 137293 -1553
rect 137411 -1671 137502 -1553
rect 137202 -1713 137502 -1671
rect 137202 -1831 137293 -1713
rect 137411 -1831 137502 -1713
rect 137202 -1842 137502 -1831
rect 139002 -2473 139302 240
rect 139002 -2591 139093 -2473
rect 139211 -2591 139302 -2473
rect 139002 -2633 139302 -2591
rect 139002 -2751 139093 -2633
rect 139211 -2751 139302 -2633
rect 139002 -2762 139302 -2751
rect 131802 -3051 131893 -2933
rect 132011 -3051 132102 -2933
rect 131802 -3093 132102 -3051
rect 131802 -3211 131893 -3093
rect 132011 -3211 132102 -3093
rect 131802 -3682 132102 -3211
rect 140802 -3393 141102 240
rect 144402 -173 144702 240
rect 144402 -291 144493 -173
rect 144611 -291 144702 -173
rect 144402 -333 144702 -291
rect 144402 -451 144493 -333
rect 144611 -451 144702 -333
rect 144402 -922 144702 -451
rect 146202 -1093 146502 240
rect 146202 -1211 146293 -1093
rect 146411 -1211 146502 -1093
rect 146202 -1253 146502 -1211
rect 146202 -1371 146293 -1253
rect 146411 -1371 146502 -1253
rect 146202 -1842 146502 -1371
rect 148002 -2013 148302 240
rect 148002 -2131 148093 -2013
rect 148211 -2131 148302 -2013
rect 148002 -2173 148302 -2131
rect 148002 -2291 148093 -2173
rect 148211 -2291 148302 -2173
rect 148002 -2762 148302 -2291
rect 140802 -3511 140893 -3393
rect 141011 -3511 141102 -3393
rect 140802 -3553 141102 -3511
rect 140802 -3671 140893 -3553
rect 141011 -3671 141102 -3553
rect 140802 -3682 141102 -3671
rect 149802 -2933 150102 240
rect 153402 -633 153702 240
rect 153402 -751 153493 -633
rect 153611 -751 153702 -633
rect 153402 -793 153702 -751
rect 153402 -911 153493 -793
rect 153611 -911 153702 -793
rect 153402 -922 153702 -911
rect 155202 -1553 155502 240
rect 155202 -1671 155293 -1553
rect 155411 -1671 155502 -1553
rect 155202 -1713 155502 -1671
rect 155202 -1831 155293 -1713
rect 155411 -1831 155502 -1713
rect 155202 -1842 155502 -1831
rect 157002 -2473 157302 240
rect 157002 -2591 157093 -2473
rect 157211 -2591 157302 -2473
rect 157002 -2633 157302 -2591
rect 157002 -2751 157093 -2633
rect 157211 -2751 157302 -2633
rect 157002 -2762 157302 -2751
rect 149802 -3051 149893 -2933
rect 150011 -3051 150102 -2933
rect 149802 -3093 150102 -3051
rect 149802 -3211 149893 -3093
rect 150011 -3211 150102 -3093
rect 149802 -3682 150102 -3211
rect 158802 -3393 159102 240
rect 162402 -173 162702 240
rect 162402 -291 162493 -173
rect 162611 -291 162702 -173
rect 162402 -333 162702 -291
rect 162402 -451 162493 -333
rect 162611 -451 162702 -333
rect 162402 -922 162702 -451
rect 164202 -1093 164502 240
rect 164202 -1211 164293 -1093
rect 164411 -1211 164502 -1093
rect 164202 -1253 164502 -1211
rect 164202 -1371 164293 -1253
rect 164411 -1371 164502 -1253
rect 164202 -1842 164502 -1371
rect 166002 -2013 166302 240
rect 166002 -2131 166093 -2013
rect 166211 -2131 166302 -2013
rect 166002 -2173 166302 -2131
rect 166002 -2291 166093 -2173
rect 166211 -2291 166302 -2173
rect 166002 -2762 166302 -2291
rect 158802 -3511 158893 -3393
rect 159011 -3511 159102 -3393
rect 158802 -3553 159102 -3511
rect 158802 -3671 158893 -3553
rect 159011 -3671 159102 -3553
rect 158802 -3682 159102 -3671
rect 167802 -2933 168102 240
rect 171402 -633 171702 240
rect 171402 -751 171493 -633
rect 171611 -751 171702 -633
rect 171402 -793 171702 -751
rect 171402 -911 171493 -793
rect 171611 -911 171702 -793
rect 171402 -922 171702 -911
rect 173202 -1553 173502 240
rect 173202 -1671 173293 -1553
rect 173411 -1671 173502 -1553
rect 173202 -1713 173502 -1671
rect 173202 -1831 173293 -1713
rect 173411 -1831 173502 -1713
rect 173202 -1842 173502 -1831
rect 175002 -2473 175302 240
rect 175002 -2591 175093 -2473
rect 175211 -2591 175302 -2473
rect 175002 -2633 175302 -2591
rect 175002 -2751 175093 -2633
rect 175211 -2751 175302 -2633
rect 175002 -2762 175302 -2751
rect 167802 -3051 167893 -2933
rect 168011 -3051 168102 -2933
rect 167802 -3093 168102 -3051
rect 167802 -3211 167893 -3093
rect 168011 -3211 168102 -3093
rect 167802 -3682 168102 -3211
rect 176802 -3393 177102 240
rect 180402 -173 180702 240
rect 180402 -291 180493 -173
rect 180611 -291 180702 -173
rect 180402 -333 180702 -291
rect 180402 -451 180493 -333
rect 180611 -451 180702 -333
rect 180402 -922 180702 -451
rect 182202 -1093 182502 240
rect 182202 -1211 182293 -1093
rect 182411 -1211 182502 -1093
rect 182202 -1253 182502 -1211
rect 182202 -1371 182293 -1253
rect 182411 -1371 182502 -1253
rect 182202 -1842 182502 -1371
rect 184002 -2013 184302 240
rect 184002 -2131 184093 -2013
rect 184211 -2131 184302 -2013
rect 184002 -2173 184302 -2131
rect 184002 -2291 184093 -2173
rect 184211 -2291 184302 -2173
rect 184002 -2762 184302 -2291
rect 176802 -3511 176893 -3393
rect 177011 -3511 177102 -3393
rect 176802 -3553 177102 -3511
rect 176802 -3671 176893 -3553
rect 177011 -3671 177102 -3553
rect 176802 -3682 177102 -3671
rect 185802 -2933 186102 240
rect 189402 -633 189702 240
rect 189402 -751 189493 -633
rect 189611 -751 189702 -633
rect 189402 -793 189702 -751
rect 189402 -911 189493 -793
rect 189611 -911 189702 -793
rect 189402 -922 189702 -911
rect 191202 -1553 191502 240
rect 191202 -1671 191293 -1553
rect 191411 -1671 191502 -1553
rect 191202 -1713 191502 -1671
rect 191202 -1831 191293 -1713
rect 191411 -1831 191502 -1713
rect 191202 -1842 191502 -1831
rect 193002 -2473 193302 240
rect 193002 -2591 193093 -2473
rect 193211 -2591 193302 -2473
rect 193002 -2633 193302 -2591
rect 193002 -2751 193093 -2633
rect 193211 -2751 193302 -2633
rect 193002 -2762 193302 -2751
rect 185802 -3051 185893 -2933
rect 186011 -3051 186102 -2933
rect 185802 -3093 186102 -3051
rect 185802 -3211 185893 -3093
rect 186011 -3211 186102 -3093
rect 185802 -3682 186102 -3211
rect 194802 -3393 195102 240
rect 198402 -173 198702 240
rect 198402 -291 198493 -173
rect 198611 -291 198702 -173
rect 198402 -333 198702 -291
rect 198402 -451 198493 -333
rect 198611 -451 198702 -333
rect 198402 -922 198702 -451
rect 200202 -1093 200502 240
rect 200202 -1211 200293 -1093
rect 200411 -1211 200502 -1093
rect 200202 -1253 200502 -1211
rect 200202 -1371 200293 -1253
rect 200411 -1371 200502 -1253
rect 200202 -1842 200502 -1371
rect 202002 -2013 202302 240
rect 202002 -2131 202093 -2013
rect 202211 -2131 202302 -2013
rect 202002 -2173 202302 -2131
rect 202002 -2291 202093 -2173
rect 202211 -2291 202302 -2173
rect 202002 -2762 202302 -2291
rect 194802 -3511 194893 -3393
rect 195011 -3511 195102 -3393
rect 194802 -3553 195102 -3511
rect 194802 -3671 194893 -3553
rect 195011 -3671 195102 -3553
rect 194802 -3682 195102 -3671
rect 203802 -2933 204102 240
rect 207402 -633 207702 240
rect 207402 -751 207493 -633
rect 207611 -751 207702 -633
rect 207402 -793 207702 -751
rect 207402 -911 207493 -793
rect 207611 -911 207702 -793
rect 207402 -922 207702 -911
rect 209202 -1553 209502 240
rect 209202 -1671 209293 -1553
rect 209411 -1671 209502 -1553
rect 209202 -1713 209502 -1671
rect 209202 -1831 209293 -1713
rect 209411 -1831 209502 -1713
rect 209202 -1842 209502 -1831
rect 211002 -2473 211302 240
rect 211002 -2591 211093 -2473
rect 211211 -2591 211302 -2473
rect 211002 -2633 211302 -2591
rect 211002 -2751 211093 -2633
rect 211211 -2751 211302 -2633
rect 211002 -2762 211302 -2751
rect 203802 -3051 203893 -2933
rect 204011 -3051 204102 -2933
rect 203802 -3093 204102 -3051
rect 203802 -3211 203893 -3093
rect 204011 -3211 204102 -3093
rect 203802 -3682 204102 -3211
rect 212802 -3393 213102 240
rect 216402 -173 216702 240
rect 216402 -291 216493 -173
rect 216611 -291 216702 -173
rect 216402 -333 216702 -291
rect 216402 -451 216493 -333
rect 216611 -451 216702 -333
rect 216402 -922 216702 -451
rect 218202 -1093 218502 240
rect 218202 -1211 218293 -1093
rect 218411 -1211 218502 -1093
rect 218202 -1253 218502 -1211
rect 218202 -1371 218293 -1253
rect 218411 -1371 218502 -1253
rect 218202 -1842 218502 -1371
rect 220002 -2013 220302 240
rect 220002 -2131 220093 -2013
rect 220211 -2131 220302 -2013
rect 220002 -2173 220302 -2131
rect 220002 -2291 220093 -2173
rect 220211 -2291 220302 -2173
rect 220002 -2762 220302 -2291
rect 212802 -3511 212893 -3393
rect 213011 -3511 213102 -3393
rect 212802 -3553 213102 -3511
rect 212802 -3671 212893 -3553
rect 213011 -3671 213102 -3553
rect 212802 -3682 213102 -3671
rect 221802 -2933 222102 240
rect 225402 -633 225702 240
rect 225402 -751 225493 -633
rect 225611 -751 225702 -633
rect 225402 -793 225702 -751
rect 225402 -911 225493 -793
rect 225611 -911 225702 -793
rect 225402 -922 225702 -911
rect 227202 -1553 227502 240
rect 227202 -1671 227293 -1553
rect 227411 -1671 227502 -1553
rect 227202 -1713 227502 -1671
rect 227202 -1831 227293 -1713
rect 227411 -1831 227502 -1713
rect 227202 -1842 227502 -1831
rect 229002 -2473 229302 240
rect 229002 -2591 229093 -2473
rect 229211 -2591 229302 -2473
rect 229002 -2633 229302 -2591
rect 229002 -2751 229093 -2633
rect 229211 -2751 229302 -2633
rect 229002 -2762 229302 -2751
rect 221802 -3051 221893 -2933
rect 222011 -3051 222102 -2933
rect 221802 -3093 222102 -3051
rect 221802 -3211 221893 -3093
rect 222011 -3211 222102 -3093
rect 221802 -3682 222102 -3211
rect 230802 -3393 231102 240
rect 234402 -173 234702 240
rect 234402 -291 234493 -173
rect 234611 -291 234702 -173
rect 234402 -333 234702 -291
rect 234402 -451 234493 -333
rect 234611 -451 234702 -333
rect 234402 -922 234702 -451
rect 236202 -1093 236502 240
rect 236202 -1211 236293 -1093
rect 236411 -1211 236502 -1093
rect 236202 -1253 236502 -1211
rect 236202 -1371 236293 -1253
rect 236411 -1371 236502 -1253
rect 236202 -1842 236502 -1371
rect 238002 -2013 238302 240
rect 238002 -2131 238093 -2013
rect 238211 -2131 238302 -2013
rect 238002 -2173 238302 -2131
rect 238002 -2291 238093 -2173
rect 238211 -2291 238302 -2173
rect 238002 -2762 238302 -2291
rect 230802 -3511 230893 -3393
rect 231011 -3511 231102 -3393
rect 230802 -3553 231102 -3511
rect 230802 -3671 230893 -3553
rect 231011 -3671 231102 -3553
rect 230802 -3682 231102 -3671
rect 239802 -2933 240102 240
rect 243402 -633 243702 240
rect 243402 -751 243493 -633
rect 243611 -751 243702 -633
rect 243402 -793 243702 -751
rect 243402 -911 243493 -793
rect 243611 -911 243702 -793
rect 243402 -922 243702 -911
rect 245202 -1553 245502 240
rect 245202 -1671 245293 -1553
rect 245411 -1671 245502 -1553
rect 245202 -1713 245502 -1671
rect 245202 -1831 245293 -1713
rect 245411 -1831 245502 -1713
rect 245202 -1842 245502 -1831
rect 247002 -2473 247302 240
rect 247002 -2591 247093 -2473
rect 247211 -2591 247302 -2473
rect 247002 -2633 247302 -2591
rect 247002 -2751 247093 -2633
rect 247211 -2751 247302 -2633
rect 247002 -2762 247302 -2751
rect 239802 -3051 239893 -2933
rect 240011 -3051 240102 -2933
rect 239802 -3093 240102 -3051
rect 239802 -3211 239893 -3093
rect 240011 -3211 240102 -3093
rect 239802 -3682 240102 -3211
rect 248802 -3393 249102 240
rect 252402 -173 252702 240
rect 252402 -291 252493 -173
rect 252611 -291 252702 -173
rect 252402 -333 252702 -291
rect 252402 -451 252493 -333
rect 252611 -451 252702 -333
rect 252402 -922 252702 -451
rect 254202 -1093 254502 240
rect 254202 -1211 254293 -1093
rect 254411 -1211 254502 -1093
rect 254202 -1253 254502 -1211
rect 254202 -1371 254293 -1253
rect 254411 -1371 254502 -1253
rect 254202 -1842 254502 -1371
rect 256002 -2013 256302 240
rect 256002 -2131 256093 -2013
rect 256211 -2131 256302 -2013
rect 256002 -2173 256302 -2131
rect 256002 -2291 256093 -2173
rect 256211 -2291 256302 -2173
rect 256002 -2762 256302 -2291
rect 248802 -3511 248893 -3393
rect 249011 -3511 249102 -3393
rect 248802 -3553 249102 -3511
rect 248802 -3671 248893 -3553
rect 249011 -3671 249102 -3553
rect 248802 -3682 249102 -3671
rect 257802 -2933 258102 240
rect 261402 -633 261702 240
rect 261402 -751 261493 -633
rect 261611 -751 261702 -633
rect 261402 -793 261702 -751
rect 261402 -911 261493 -793
rect 261611 -911 261702 -793
rect 261402 -922 261702 -911
rect 263202 -1553 263502 240
rect 263202 -1671 263293 -1553
rect 263411 -1671 263502 -1553
rect 263202 -1713 263502 -1671
rect 263202 -1831 263293 -1713
rect 263411 -1831 263502 -1713
rect 263202 -1842 263502 -1831
rect 265002 -2473 265302 240
rect 265002 -2591 265093 -2473
rect 265211 -2591 265302 -2473
rect 265002 -2633 265302 -2591
rect 265002 -2751 265093 -2633
rect 265211 -2751 265302 -2633
rect 265002 -2762 265302 -2751
rect 257802 -3051 257893 -2933
rect 258011 -3051 258102 -2933
rect 257802 -3093 258102 -3051
rect 257802 -3211 257893 -3093
rect 258011 -3211 258102 -3093
rect 257802 -3682 258102 -3211
rect 266802 -3393 267102 240
rect 270402 -173 270702 240
rect 270402 -291 270493 -173
rect 270611 -291 270702 -173
rect 270402 -333 270702 -291
rect 270402 -451 270493 -333
rect 270611 -451 270702 -333
rect 270402 -922 270702 -451
rect 272202 -1093 272502 240
rect 272202 -1211 272293 -1093
rect 272411 -1211 272502 -1093
rect 272202 -1253 272502 -1211
rect 272202 -1371 272293 -1253
rect 272411 -1371 272502 -1253
rect 272202 -1842 272502 -1371
rect 274002 -2013 274302 240
rect 274002 -2131 274093 -2013
rect 274211 -2131 274302 -2013
rect 274002 -2173 274302 -2131
rect 274002 -2291 274093 -2173
rect 274211 -2291 274302 -2173
rect 274002 -2762 274302 -2291
rect 266802 -3511 266893 -3393
rect 267011 -3511 267102 -3393
rect 266802 -3553 267102 -3511
rect 266802 -3671 266893 -3553
rect 267011 -3671 267102 -3553
rect 266802 -3682 267102 -3671
rect 275802 -2933 276102 240
rect 279402 -633 279702 240
rect 279402 -751 279493 -633
rect 279611 -751 279702 -633
rect 279402 -793 279702 -751
rect 279402 -911 279493 -793
rect 279611 -911 279702 -793
rect 279402 -922 279702 -911
rect 281202 -1553 281502 240
rect 281202 -1671 281293 -1553
rect 281411 -1671 281502 -1553
rect 281202 -1713 281502 -1671
rect 281202 -1831 281293 -1713
rect 281411 -1831 281502 -1713
rect 281202 -1842 281502 -1831
rect 283002 -2473 283302 240
rect 283002 -2591 283093 -2473
rect 283211 -2591 283302 -2473
rect 283002 -2633 283302 -2591
rect 283002 -2751 283093 -2633
rect 283211 -2751 283302 -2633
rect 283002 -2762 283302 -2751
rect 275802 -3051 275893 -2933
rect 276011 -3051 276102 -2933
rect 275802 -3093 276102 -3051
rect 275802 -3211 275893 -3093
rect 276011 -3211 276102 -3093
rect 275802 -3682 276102 -3211
rect 284802 -3393 285102 240
rect 288402 -173 288702 240
rect 288402 -291 288493 -173
rect 288611 -291 288702 -173
rect 288402 -333 288702 -291
rect 288402 -451 288493 -333
rect 288611 -451 288702 -333
rect 288402 -922 288702 -451
rect 290202 -1093 290502 240
rect 292660 -173 292960 949
rect 292660 -291 292751 -173
rect 292869 -291 292960 -173
rect 292660 -333 292960 -291
rect 292660 -451 292751 -333
rect 292869 -451 292960 -333
rect 292660 -462 292960 -451
rect 293120 334227 293420 352601
rect 293120 334109 293211 334227
rect 293329 334109 293420 334227
rect 293120 334067 293420 334109
rect 293120 333949 293211 334067
rect 293329 333949 293420 334067
rect 293120 316227 293420 333949
rect 293120 316109 293211 316227
rect 293329 316109 293420 316227
rect 293120 316067 293420 316109
rect 293120 315949 293211 316067
rect 293329 315949 293420 316067
rect 293120 298227 293420 315949
rect 293120 298109 293211 298227
rect 293329 298109 293420 298227
rect 293120 298067 293420 298109
rect 293120 297949 293211 298067
rect 293329 297949 293420 298067
rect 293120 280227 293420 297949
rect 293120 280109 293211 280227
rect 293329 280109 293420 280227
rect 293120 280067 293420 280109
rect 293120 279949 293211 280067
rect 293329 279949 293420 280067
rect 293120 262227 293420 279949
rect 293120 262109 293211 262227
rect 293329 262109 293420 262227
rect 293120 262067 293420 262109
rect 293120 261949 293211 262067
rect 293329 261949 293420 262067
rect 293120 244227 293420 261949
rect 293120 244109 293211 244227
rect 293329 244109 293420 244227
rect 293120 244067 293420 244109
rect 293120 243949 293211 244067
rect 293329 243949 293420 244067
rect 293120 226227 293420 243949
rect 293120 226109 293211 226227
rect 293329 226109 293420 226227
rect 293120 226067 293420 226109
rect 293120 225949 293211 226067
rect 293329 225949 293420 226067
rect 293120 208227 293420 225949
rect 293120 208109 293211 208227
rect 293329 208109 293420 208227
rect 293120 208067 293420 208109
rect 293120 207949 293211 208067
rect 293329 207949 293420 208067
rect 293120 190227 293420 207949
rect 293120 190109 293211 190227
rect 293329 190109 293420 190227
rect 293120 190067 293420 190109
rect 293120 189949 293211 190067
rect 293329 189949 293420 190067
rect 293120 172227 293420 189949
rect 293120 172109 293211 172227
rect 293329 172109 293420 172227
rect 293120 172067 293420 172109
rect 293120 171949 293211 172067
rect 293329 171949 293420 172067
rect 293120 154227 293420 171949
rect 293120 154109 293211 154227
rect 293329 154109 293420 154227
rect 293120 154067 293420 154109
rect 293120 153949 293211 154067
rect 293329 153949 293420 154067
rect 293120 136227 293420 153949
rect 293120 136109 293211 136227
rect 293329 136109 293420 136227
rect 293120 136067 293420 136109
rect 293120 135949 293211 136067
rect 293329 135949 293420 136067
rect 293120 118227 293420 135949
rect 293120 118109 293211 118227
rect 293329 118109 293420 118227
rect 293120 118067 293420 118109
rect 293120 117949 293211 118067
rect 293329 117949 293420 118067
rect 293120 100227 293420 117949
rect 293120 100109 293211 100227
rect 293329 100109 293420 100227
rect 293120 100067 293420 100109
rect 293120 99949 293211 100067
rect 293329 99949 293420 100067
rect 293120 82227 293420 99949
rect 293120 82109 293211 82227
rect 293329 82109 293420 82227
rect 293120 82067 293420 82109
rect 293120 81949 293211 82067
rect 293329 81949 293420 82067
rect 293120 64227 293420 81949
rect 293120 64109 293211 64227
rect 293329 64109 293420 64227
rect 293120 64067 293420 64109
rect 293120 63949 293211 64067
rect 293329 63949 293420 64067
rect 293120 46227 293420 63949
rect 293120 46109 293211 46227
rect 293329 46109 293420 46227
rect 293120 46067 293420 46109
rect 293120 45949 293211 46067
rect 293329 45949 293420 46067
rect 293120 28227 293420 45949
rect 293120 28109 293211 28227
rect 293329 28109 293420 28227
rect 293120 28067 293420 28109
rect 293120 27949 293211 28067
rect 293329 27949 293420 28067
rect 293120 10227 293420 27949
rect 293120 10109 293211 10227
rect 293329 10109 293420 10227
rect 293120 10067 293420 10109
rect 293120 9949 293211 10067
rect 293329 9949 293420 10067
rect 293120 -633 293420 9949
rect 293120 -751 293211 -633
rect 293329 -751 293420 -633
rect 293120 -793 293420 -751
rect 293120 -911 293211 -793
rect 293329 -911 293420 -793
rect 293120 -922 293420 -911
rect 293580 345027 293880 353061
rect 293580 344909 293671 345027
rect 293789 344909 293880 345027
rect 293580 344867 293880 344909
rect 293580 344749 293671 344867
rect 293789 344749 293880 344867
rect 293580 327027 293880 344749
rect 293580 326909 293671 327027
rect 293789 326909 293880 327027
rect 293580 326867 293880 326909
rect 293580 326749 293671 326867
rect 293789 326749 293880 326867
rect 293580 309027 293880 326749
rect 293580 308909 293671 309027
rect 293789 308909 293880 309027
rect 293580 308867 293880 308909
rect 293580 308749 293671 308867
rect 293789 308749 293880 308867
rect 293580 291027 293880 308749
rect 293580 290909 293671 291027
rect 293789 290909 293880 291027
rect 293580 290867 293880 290909
rect 293580 290749 293671 290867
rect 293789 290749 293880 290867
rect 293580 273027 293880 290749
rect 293580 272909 293671 273027
rect 293789 272909 293880 273027
rect 293580 272867 293880 272909
rect 293580 272749 293671 272867
rect 293789 272749 293880 272867
rect 293580 255027 293880 272749
rect 293580 254909 293671 255027
rect 293789 254909 293880 255027
rect 293580 254867 293880 254909
rect 293580 254749 293671 254867
rect 293789 254749 293880 254867
rect 293580 237027 293880 254749
rect 293580 236909 293671 237027
rect 293789 236909 293880 237027
rect 293580 236867 293880 236909
rect 293580 236749 293671 236867
rect 293789 236749 293880 236867
rect 293580 219027 293880 236749
rect 293580 218909 293671 219027
rect 293789 218909 293880 219027
rect 293580 218867 293880 218909
rect 293580 218749 293671 218867
rect 293789 218749 293880 218867
rect 293580 201027 293880 218749
rect 293580 200909 293671 201027
rect 293789 200909 293880 201027
rect 293580 200867 293880 200909
rect 293580 200749 293671 200867
rect 293789 200749 293880 200867
rect 293580 183027 293880 200749
rect 293580 182909 293671 183027
rect 293789 182909 293880 183027
rect 293580 182867 293880 182909
rect 293580 182749 293671 182867
rect 293789 182749 293880 182867
rect 293580 165027 293880 182749
rect 293580 164909 293671 165027
rect 293789 164909 293880 165027
rect 293580 164867 293880 164909
rect 293580 164749 293671 164867
rect 293789 164749 293880 164867
rect 293580 147027 293880 164749
rect 293580 146909 293671 147027
rect 293789 146909 293880 147027
rect 293580 146867 293880 146909
rect 293580 146749 293671 146867
rect 293789 146749 293880 146867
rect 293580 129027 293880 146749
rect 293580 128909 293671 129027
rect 293789 128909 293880 129027
rect 293580 128867 293880 128909
rect 293580 128749 293671 128867
rect 293789 128749 293880 128867
rect 293580 111027 293880 128749
rect 293580 110909 293671 111027
rect 293789 110909 293880 111027
rect 293580 110867 293880 110909
rect 293580 110749 293671 110867
rect 293789 110749 293880 110867
rect 293580 93027 293880 110749
rect 293580 92909 293671 93027
rect 293789 92909 293880 93027
rect 293580 92867 293880 92909
rect 293580 92749 293671 92867
rect 293789 92749 293880 92867
rect 293580 75027 293880 92749
rect 293580 74909 293671 75027
rect 293789 74909 293880 75027
rect 293580 74867 293880 74909
rect 293580 74749 293671 74867
rect 293789 74749 293880 74867
rect 293580 57027 293880 74749
rect 293580 56909 293671 57027
rect 293789 56909 293880 57027
rect 293580 56867 293880 56909
rect 293580 56749 293671 56867
rect 293789 56749 293880 56867
rect 293580 39027 293880 56749
rect 293580 38909 293671 39027
rect 293789 38909 293880 39027
rect 293580 38867 293880 38909
rect 293580 38749 293671 38867
rect 293789 38749 293880 38867
rect 293580 21027 293880 38749
rect 293580 20909 293671 21027
rect 293789 20909 293880 21027
rect 293580 20867 293880 20909
rect 293580 20749 293671 20867
rect 293789 20749 293880 20867
rect 293580 3027 293880 20749
rect 293580 2909 293671 3027
rect 293789 2909 293880 3027
rect 293580 2867 293880 2909
rect 293580 2749 293671 2867
rect 293789 2749 293880 2867
rect 290202 -1211 290293 -1093
rect 290411 -1211 290502 -1093
rect 290202 -1253 290502 -1211
rect 290202 -1371 290293 -1253
rect 290411 -1371 290502 -1253
rect 290202 -1842 290502 -1371
rect 293580 -1093 293880 2749
rect 293580 -1211 293671 -1093
rect 293789 -1211 293880 -1093
rect 293580 -1253 293880 -1211
rect 293580 -1371 293671 -1253
rect 293789 -1371 293880 -1253
rect 293580 -1382 293880 -1371
rect 294040 336027 294340 353521
rect 294040 335909 294131 336027
rect 294249 335909 294340 336027
rect 294040 335867 294340 335909
rect 294040 335749 294131 335867
rect 294249 335749 294340 335867
rect 294040 318027 294340 335749
rect 294040 317909 294131 318027
rect 294249 317909 294340 318027
rect 294040 317867 294340 317909
rect 294040 317749 294131 317867
rect 294249 317749 294340 317867
rect 294040 300027 294340 317749
rect 294040 299909 294131 300027
rect 294249 299909 294340 300027
rect 294040 299867 294340 299909
rect 294040 299749 294131 299867
rect 294249 299749 294340 299867
rect 294040 282027 294340 299749
rect 294040 281909 294131 282027
rect 294249 281909 294340 282027
rect 294040 281867 294340 281909
rect 294040 281749 294131 281867
rect 294249 281749 294340 281867
rect 294040 264027 294340 281749
rect 294040 263909 294131 264027
rect 294249 263909 294340 264027
rect 294040 263867 294340 263909
rect 294040 263749 294131 263867
rect 294249 263749 294340 263867
rect 294040 246027 294340 263749
rect 294040 245909 294131 246027
rect 294249 245909 294340 246027
rect 294040 245867 294340 245909
rect 294040 245749 294131 245867
rect 294249 245749 294340 245867
rect 294040 228027 294340 245749
rect 294040 227909 294131 228027
rect 294249 227909 294340 228027
rect 294040 227867 294340 227909
rect 294040 227749 294131 227867
rect 294249 227749 294340 227867
rect 294040 210027 294340 227749
rect 294040 209909 294131 210027
rect 294249 209909 294340 210027
rect 294040 209867 294340 209909
rect 294040 209749 294131 209867
rect 294249 209749 294340 209867
rect 294040 192027 294340 209749
rect 294040 191909 294131 192027
rect 294249 191909 294340 192027
rect 294040 191867 294340 191909
rect 294040 191749 294131 191867
rect 294249 191749 294340 191867
rect 294040 174027 294340 191749
rect 294040 173909 294131 174027
rect 294249 173909 294340 174027
rect 294040 173867 294340 173909
rect 294040 173749 294131 173867
rect 294249 173749 294340 173867
rect 294040 156027 294340 173749
rect 294040 155909 294131 156027
rect 294249 155909 294340 156027
rect 294040 155867 294340 155909
rect 294040 155749 294131 155867
rect 294249 155749 294340 155867
rect 294040 138027 294340 155749
rect 294040 137909 294131 138027
rect 294249 137909 294340 138027
rect 294040 137867 294340 137909
rect 294040 137749 294131 137867
rect 294249 137749 294340 137867
rect 294040 120027 294340 137749
rect 294040 119909 294131 120027
rect 294249 119909 294340 120027
rect 294040 119867 294340 119909
rect 294040 119749 294131 119867
rect 294249 119749 294340 119867
rect 294040 102027 294340 119749
rect 294040 101909 294131 102027
rect 294249 101909 294340 102027
rect 294040 101867 294340 101909
rect 294040 101749 294131 101867
rect 294249 101749 294340 101867
rect 294040 84027 294340 101749
rect 294040 83909 294131 84027
rect 294249 83909 294340 84027
rect 294040 83867 294340 83909
rect 294040 83749 294131 83867
rect 294249 83749 294340 83867
rect 294040 66027 294340 83749
rect 294040 65909 294131 66027
rect 294249 65909 294340 66027
rect 294040 65867 294340 65909
rect 294040 65749 294131 65867
rect 294249 65749 294340 65867
rect 294040 48027 294340 65749
rect 294040 47909 294131 48027
rect 294249 47909 294340 48027
rect 294040 47867 294340 47909
rect 294040 47749 294131 47867
rect 294249 47749 294340 47867
rect 294040 30027 294340 47749
rect 294040 29909 294131 30027
rect 294249 29909 294340 30027
rect 294040 29867 294340 29909
rect 294040 29749 294131 29867
rect 294249 29749 294340 29867
rect 294040 12027 294340 29749
rect 294040 11909 294131 12027
rect 294249 11909 294340 12027
rect 294040 11867 294340 11909
rect 294040 11749 294131 11867
rect 294249 11749 294340 11867
rect 294040 -1553 294340 11749
rect 294040 -1671 294131 -1553
rect 294249 -1671 294340 -1553
rect 294040 -1713 294340 -1671
rect 294040 -1831 294131 -1713
rect 294249 -1831 294340 -1713
rect 294040 -1842 294340 -1831
rect 294500 346827 294800 353981
rect 294500 346709 294591 346827
rect 294709 346709 294800 346827
rect 294500 346667 294800 346709
rect 294500 346549 294591 346667
rect 294709 346549 294800 346667
rect 294500 328827 294800 346549
rect 294500 328709 294591 328827
rect 294709 328709 294800 328827
rect 294500 328667 294800 328709
rect 294500 328549 294591 328667
rect 294709 328549 294800 328667
rect 294500 310827 294800 328549
rect 294500 310709 294591 310827
rect 294709 310709 294800 310827
rect 294500 310667 294800 310709
rect 294500 310549 294591 310667
rect 294709 310549 294800 310667
rect 294500 292827 294800 310549
rect 294500 292709 294591 292827
rect 294709 292709 294800 292827
rect 294500 292667 294800 292709
rect 294500 292549 294591 292667
rect 294709 292549 294800 292667
rect 294500 274827 294800 292549
rect 294500 274709 294591 274827
rect 294709 274709 294800 274827
rect 294500 274667 294800 274709
rect 294500 274549 294591 274667
rect 294709 274549 294800 274667
rect 294500 256827 294800 274549
rect 294500 256709 294591 256827
rect 294709 256709 294800 256827
rect 294500 256667 294800 256709
rect 294500 256549 294591 256667
rect 294709 256549 294800 256667
rect 294500 238827 294800 256549
rect 294500 238709 294591 238827
rect 294709 238709 294800 238827
rect 294500 238667 294800 238709
rect 294500 238549 294591 238667
rect 294709 238549 294800 238667
rect 294500 220827 294800 238549
rect 294500 220709 294591 220827
rect 294709 220709 294800 220827
rect 294500 220667 294800 220709
rect 294500 220549 294591 220667
rect 294709 220549 294800 220667
rect 294500 202827 294800 220549
rect 294500 202709 294591 202827
rect 294709 202709 294800 202827
rect 294500 202667 294800 202709
rect 294500 202549 294591 202667
rect 294709 202549 294800 202667
rect 294500 184827 294800 202549
rect 294500 184709 294591 184827
rect 294709 184709 294800 184827
rect 294500 184667 294800 184709
rect 294500 184549 294591 184667
rect 294709 184549 294800 184667
rect 294500 166827 294800 184549
rect 294500 166709 294591 166827
rect 294709 166709 294800 166827
rect 294500 166667 294800 166709
rect 294500 166549 294591 166667
rect 294709 166549 294800 166667
rect 294500 148827 294800 166549
rect 294500 148709 294591 148827
rect 294709 148709 294800 148827
rect 294500 148667 294800 148709
rect 294500 148549 294591 148667
rect 294709 148549 294800 148667
rect 294500 130827 294800 148549
rect 294500 130709 294591 130827
rect 294709 130709 294800 130827
rect 294500 130667 294800 130709
rect 294500 130549 294591 130667
rect 294709 130549 294800 130667
rect 294500 112827 294800 130549
rect 294500 112709 294591 112827
rect 294709 112709 294800 112827
rect 294500 112667 294800 112709
rect 294500 112549 294591 112667
rect 294709 112549 294800 112667
rect 294500 94827 294800 112549
rect 294500 94709 294591 94827
rect 294709 94709 294800 94827
rect 294500 94667 294800 94709
rect 294500 94549 294591 94667
rect 294709 94549 294800 94667
rect 294500 76827 294800 94549
rect 294500 76709 294591 76827
rect 294709 76709 294800 76827
rect 294500 76667 294800 76709
rect 294500 76549 294591 76667
rect 294709 76549 294800 76667
rect 294500 58827 294800 76549
rect 294500 58709 294591 58827
rect 294709 58709 294800 58827
rect 294500 58667 294800 58709
rect 294500 58549 294591 58667
rect 294709 58549 294800 58667
rect 294500 40827 294800 58549
rect 294500 40709 294591 40827
rect 294709 40709 294800 40827
rect 294500 40667 294800 40709
rect 294500 40549 294591 40667
rect 294709 40549 294800 40667
rect 294500 22827 294800 40549
rect 294500 22709 294591 22827
rect 294709 22709 294800 22827
rect 294500 22667 294800 22709
rect 294500 22549 294591 22667
rect 294709 22549 294800 22667
rect 294500 4827 294800 22549
rect 294500 4709 294591 4827
rect 294709 4709 294800 4827
rect 294500 4667 294800 4709
rect 294500 4549 294591 4667
rect 294709 4549 294800 4667
rect 294500 -2013 294800 4549
rect 294500 -2131 294591 -2013
rect 294709 -2131 294800 -2013
rect 294500 -2173 294800 -2131
rect 294500 -2291 294591 -2173
rect 294709 -2291 294800 -2173
rect 294500 -2302 294800 -2291
rect 294960 337827 295260 354441
rect 294960 337709 295051 337827
rect 295169 337709 295260 337827
rect 294960 337667 295260 337709
rect 294960 337549 295051 337667
rect 295169 337549 295260 337667
rect 294960 319827 295260 337549
rect 294960 319709 295051 319827
rect 295169 319709 295260 319827
rect 294960 319667 295260 319709
rect 294960 319549 295051 319667
rect 295169 319549 295260 319667
rect 294960 301827 295260 319549
rect 294960 301709 295051 301827
rect 295169 301709 295260 301827
rect 294960 301667 295260 301709
rect 294960 301549 295051 301667
rect 295169 301549 295260 301667
rect 294960 283827 295260 301549
rect 294960 283709 295051 283827
rect 295169 283709 295260 283827
rect 294960 283667 295260 283709
rect 294960 283549 295051 283667
rect 295169 283549 295260 283667
rect 294960 265827 295260 283549
rect 294960 265709 295051 265827
rect 295169 265709 295260 265827
rect 294960 265667 295260 265709
rect 294960 265549 295051 265667
rect 295169 265549 295260 265667
rect 294960 247827 295260 265549
rect 294960 247709 295051 247827
rect 295169 247709 295260 247827
rect 294960 247667 295260 247709
rect 294960 247549 295051 247667
rect 295169 247549 295260 247667
rect 294960 229827 295260 247549
rect 294960 229709 295051 229827
rect 295169 229709 295260 229827
rect 294960 229667 295260 229709
rect 294960 229549 295051 229667
rect 295169 229549 295260 229667
rect 294960 211827 295260 229549
rect 294960 211709 295051 211827
rect 295169 211709 295260 211827
rect 294960 211667 295260 211709
rect 294960 211549 295051 211667
rect 295169 211549 295260 211667
rect 294960 193827 295260 211549
rect 294960 193709 295051 193827
rect 295169 193709 295260 193827
rect 294960 193667 295260 193709
rect 294960 193549 295051 193667
rect 295169 193549 295260 193667
rect 294960 175827 295260 193549
rect 294960 175709 295051 175827
rect 295169 175709 295260 175827
rect 294960 175667 295260 175709
rect 294960 175549 295051 175667
rect 295169 175549 295260 175667
rect 294960 157827 295260 175549
rect 294960 157709 295051 157827
rect 295169 157709 295260 157827
rect 294960 157667 295260 157709
rect 294960 157549 295051 157667
rect 295169 157549 295260 157667
rect 294960 139827 295260 157549
rect 294960 139709 295051 139827
rect 295169 139709 295260 139827
rect 294960 139667 295260 139709
rect 294960 139549 295051 139667
rect 295169 139549 295260 139667
rect 294960 121827 295260 139549
rect 294960 121709 295051 121827
rect 295169 121709 295260 121827
rect 294960 121667 295260 121709
rect 294960 121549 295051 121667
rect 295169 121549 295260 121667
rect 294960 103827 295260 121549
rect 294960 103709 295051 103827
rect 295169 103709 295260 103827
rect 294960 103667 295260 103709
rect 294960 103549 295051 103667
rect 295169 103549 295260 103667
rect 294960 85827 295260 103549
rect 294960 85709 295051 85827
rect 295169 85709 295260 85827
rect 294960 85667 295260 85709
rect 294960 85549 295051 85667
rect 295169 85549 295260 85667
rect 294960 67827 295260 85549
rect 294960 67709 295051 67827
rect 295169 67709 295260 67827
rect 294960 67667 295260 67709
rect 294960 67549 295051 67667
rect 295169 67549 295260 67667
rect 294960 49827 295260 67549
rect 294960 49709 295051 49827
rect 295169 49709 295260 49827
rect 294960 49667 295260 49709
rect 294960 49549 295051 49667
rect 295169 49549 295260 49667
rect 294960 31827 295260 49549
rect 294960 31709 295051 31827
rect 295169 31709 295260 31827
rect 294960 31667 295260 31709
rect 294960 31549 295051 31667
rect 295169 31549 295260 31667
rect 294960 13827 295260 31549
rect 294960 13709 295051 13827
rect 295169 13709 295260 13827
rect 294960 13667 295260 13709
rect 294960 13549 295051 13667
rect 295169 13549 295260 13667
rect 294960 -2473 295260 13549
rect 294960 -2591 295051 -2473
rect 295169 -2591 295260 -2473
rect 294960 -2633 295260 -2591
rect 294960 -2751 295051 -2633
rect 295169 -2751 295260 -2633
rect 294960 -2762 295260 -2751
rect 295420 348627 295720 354901
rect 295420 348509 295511 348627
rect 295629 348509 295720 348627
rect 295420 348467 295720 348509
rect 295420 348349 295511 348467
rect 295629 348349 295720 348467
rect 295420 330627 295720 348349
rect 295420 330509 295511 330627
rect 295629 330509 295720 330627
rect 295420 330467 295720 330509
rect 295420 330349 295511 330467
rect 295629 330349 295720 330467
rect 295420 312627 295720 330349
rect 295420 312509 295511 312627
rect 295629 312509 295720 312627
rect 295420 312467 295720 312509
rect 295420 312349 295511 312467
rect 295629 312349 295720 312467
rect 295420 294627 295720 312349
rect 295420 294509 295511 294627
rect 295629 294509 295720 294627
rect 295420 294467 295720 294509
rect 295420 294349 295511 294467
rect 295629 294349 295720 294467
rect 295420 276627 295720 294349
rect 295420 276509 295511 276627
rect 295629 276509 295720 276627
rect 295420 276467 295720 276509
rect 295420 276349 295511 276467
rect 295629 276349 295720 276467
rect 295420 258627 295720 276349
rect 295420 258509 295511 258627
rect 295629 258509 295720 258627
rect 295420 258467 295720 258509
rect 295420 258349 295511 258467
rect 295629 258349 295720 258467
rect 295420 240627 295720 258349
rect 295420 240509 295511 240627
rect 295629 240509 295720 240627
rect 295420 240467 295720 240509
rect 295420 240349 295511 240467
rect 295629 240349 295720 240467
rect 295420 222627 295720 240349
rect 295420 222509 295511 222627
rect 295629 222509 295720 222627
rect 295420 222467 295720 222509
rect 295420 222349 295511 222467
rect 295629 222349 295720 222467
rect 295420 204627 295720 222349
rect 295420 204509 295511 204627
rect 295629 204509 295720 204627
rect 295420 204467 295720 204509
rect 295420 204349 295511 204467
rect 295629 204349 295720 204467
rect 295420 186627 295720 204349
rect 295420 186509 295511 186627
rect 295629 186509 295720 186627
rect 295420 186467 295720 186509
rect 295420 186349 295511 186467
rect 295629 186349 295720 186467
rect 295420 168627 295720 186349
rect 295420 168509 295511 168627
rect 295629 168509 295720 168627
rect 295420 168467 295720 168509
rect 295420 168349 295511 168467
rect 295629 168349 295720 168467
rect 295420 150627 295720 168349
rect 295420 150509 295511 150627
rect 295629 150509 295720 150627
rect 295420 150467 295720 150509
rect 295420 150349 295511 150467
rect 295629 150349 295720 150467
rect 295420 132627 295720 150349
rect 295420 132509 295511 132627
rect 295629 132509 295720 132627
rect 295420 132467 295720 132509
rect 295420 132349 295511 132467
rect 295629 132349 295720 132467
rect 295420 114627 295720 132349
rect 295420 114509 295511 114627
rect 295629 114509 295720 114627
rect 295420 114467 295720 114509
rect 295420 114349 295511 114467
rect 295629 114349 295720 114467
rect 295420 96627 295720 114349
rect 295420 96509 295511 96627
rect 295629 96509 295720 96627
rect 295420 96467 295720 96509
rect 295420 96349 295511 96467
rect 295629 96349 295720 96467
rect 295420 78627 295720 96349
rect 295420 78509 295511 78627
rect 295629 78509 295720 78627
rect 295420 78467 295720 78509
rect 295420 78349 295511 78467
rect 295629 78349 295720 78467
rect 295420 60627 295720 78349
rect 295420 60509 295511 60627
rect 295629 60509 295720 60627
rect 295420 60467 295720 60509
rect 295420 60349 295511 60467
rect 295629 60349 295720 60467
rect 295420 42627 295720 60349
rect 295420 42509 295511 42627
rect 295629 42509 295720 42627
rect 295420 42467 295720 42509
rect 295420 42349 295511 42467
rect 295629 42349 295720 42467
rect 295420 24627 295720 42349
rect 295420 24509 295511 24627
rect 295629 24509 295720 24627
rect 295420 24467 295720 24509
rect 295420 24349 295511 24467
rect 295629 24349 295720 24467
rect 295420 6627 295720 24349
rect 295420 6509 295511 6627
rect 295629 6509 295720 6627
rect 295420 6467 295720 6509
rect 295420 6349 295511 6467
rect 295629 6349 295720 6467
rect 295420 -2933 295720 6349
rect 295420 -3051 295511 -2933
rect 295629 -3051 295720 -2933
rect 295420 -3093 295720 -3051
rect 295420 -3211 295511 -3093
rect 295629 -3211 295720 -3093
rect 295420 -3222 295720 -3211
rect 295880 339627 296180 355361
rect 295880 339509 295971 339627
rect 296089 339509 296180 339627
rect 295880 339467 296180 339509
rect 295880 339349 295971 339467
rect 296089 339349 296180 339467
rect 295880 321627 296180 339349
rect 295880 321509 295971 321627
rect 296089 321509 296180 321627
rect 295880 321467 296180 321509
rect 295880 321349 295971 321467
rect 296089 321349 296180 321467
rect 295880 303627 296180 321349
rect 295880 303509 295971 303627
rect 296089 303509 296180 303627
rect 295880 303467 296180 303509
rect 295880 303349 295971 303467
rect 296089 303349 296180 303467
rect 295880 285627 296180 303349
rect 295880 285509 295971 285627
rect 296089 285509 296180 285627
rect 295880 285467 296180 285509
rect 295880 285349 295971 285467
rect 296089 285349 296180 285467
rect 295880 267627 296180 285349
rect 295880 267509 295971 267627
rect 296089 267509 296180 267627
rect 295880 267467 296180 267509
rect 295880 267349 295971 267467
rect 296089 267349 296180 267467
rect 295880 249627 296180 267349
rect 295880 249509 295971 249627
rect 296089 249509 296180 249627
rect 295880 249467 296180 249509
rect 295880 249349 295971 249467
rect 296089 249349 296180 249467
rect 295880 231627 296180 249349
rect 295880 231509 295971 231627
rect 296089 231509 296180 231627
rect 295880 231467 296180 231509
rect 295880 231349 295971 231467
rect 296089 231349 296180 231467
rect 295880 213627 296180 231349
rect 295880 213509 295971 213627
rect 296089 213509 296180 213627
rect 295880 213467 296180 213509
rect 295880 213349 295971 213467
rect 296089 213349 296180 213467
rect 295880 195627 296180 213349
rect 295880 195509 295971 195627
rect 296089 195509 296180 195627
rect 295880 195467 296180 195509
rect 295880 195349 295971 195467
rect 296089 195349 296180 195467
rect 295880 177627 296180 195349
rect 295880 177509 295971 177627
rect 296089 177509 296180 177627
rect 295880 177467 296180 177509
rect 295880 177349 295971 177467
rect 296089 177349 296180 177467
rect 295880 159627 296180 177349
rect 295880 159509 295971 159627
rect 296089 159509 296180 159627
rect 295880 159467 296180 159509
rect 295880 159349 295971 159467
rect 296089 159349 296180 159467
rect 295880 141627 296180 159349
rect 295880 141509 295971 141627
rect 296089 141509 296180 141627
rect 295880 141467 296180 141509
rect 295880 141349 295971 141467
rect 296089 141349 296180 141467
rect 295880 123627 296180 141349
rect 295880 123509 295971 123627
rect 296089 123509 296180 123627
rect 295880 123467 296180 123509
rect 295880 123349 295971 123467
rect 296089 123349 296180 123467
rect 295880 105627 296180 123349
rect 295880 105509 295971 105627
rect 296089 105509 296180 105627
rect 295880 105467 296180 105509
rect 295880 105349 295971 105467
rect 296089 105349 296180 105467
rect 295880 87627 296180 105349
rect 295880 87509 295971 87627
rect 296089 87509 296180 87627
rect 295880 87467 296180 87509
rect 295880 87349 295971 87467
rect 296089 87349 296180 87467
rect 295880 69627 296180 87349
rect 295880 69509 295971 69627
rect 296089 69509 296180 69627
rect 295880 69467 296180 69509
rect 295880 69349 295971 69467
rect 296089 69349 296180 69467
rect 295880 51627 296180 69349
rect 295880 51509 295971 51627
rect 296089 51509 296180 51627
rect 295880 51467 296180 51509
rect 295880 51349 295971 51467
rect 296089 51349 296180 51467
rect 295880 33627 296180 51349
rect 295880 33509 295971 33627
rect 296089 33509 296180 33627
rect 295880 33467 296180 33509
rect 295880 33349 295971 33467
rect 296089 33349 296180 33467
rect 295880 15627 296180 33349
rect 295880 15509 295971 15627
rect 296089 15509 296180 15627
rect 295880 15467 296180 15509
rect 295880 15349 295971 15467
rect 296089 15349 296180 15467
rect 284802 -3511 284893 -3393
rect 285011 -3511 285102 -3393
rect 284802 -3553 285102 -3511
rect 284802 -3671 284893 -3553
rect 285011 -3671 285102 -3553
rect 284802 -3682 285102 -3671
rect 295880 -3393 296180 15349
rect 295880 -3511 295971 -3393
rect 296089 -3511 296180 -3393
rect 295880 -3553 296180 -3511
rect 295880 -3671 295971 -3553
rect 296089 -3671 296180 -3553
rect 295880 -3682 296180 -3671
<< via4 >>
rect -4127 355521 -4009 355639
rect -4127 355361 -4009 355479
rect -4127 339509 -4009 339627
rect -4127 339349 -4009 339467
rect -4127 321509 -4009 321627
rect -4127 321349 -4009 321467
rect -4127 303509 -4009 303627
rect -4127 303349 -4009 303467
rect -4127 285509 -4009 285627
rect -4127 285349 -4009 285467
rect -4127 267509 -4009 267627
rect -4127 267349 -4009 267467
rect -4127 249509 -4009 249627
rect -4127 249349 -4009 249467
rect -4127 231509 -4009 231627
rect -4127 231349 -4009 231467
rect -4127 213509 -4009 213627
rect -4127 213349 -4009 213467
rect -4127 195509 -4009 195627
rect -4127 195349 -4009 195467
rect -4127 177509 -4009 177627
rect -4127 177349 -4009 177467
rect -4127 159509 -4009 159627
rect -4127 159349 -4009 159467
rect -4127 141509 -4009 141627
rect -4127 141349 -4009 141467
rect -4127 123509 -4009 123627
rect -4127 123349 -4009 123467
rect -4127 105509 -4009 105627
rect -4127 105349 -4009 105467
rect -4127 87509 -4009 87627
rect -4127 87349 -4009 87467
rect -4127 69509 -4009 69627
rect -4127 69349 -4009 69467
rect -4127 51509 -4009 51627
rect -4127 51349 -4009 51467
rect -4127 33509 -4009 33627
rect -4127 33349 -4009 33467
rect -4127 15509 -4009 15627
rect -4127 15349 -4009 15467
rect -3667 355061 -3549 355179
rect -3667 354901 -3549 355019
rect 5893 355061 6011 355179
rect 5893 354901 6011 355019
rect -3667 348509 -3549 348627
rect -3667 348349 -3549 348467
rect -3667 330509 -3549 330627
rect -3667 330349 -3549 330467
rect -3667 312509 -3549 312627
rect -3667 312349 -3549 312467
rect -3667 294509 -3549 294627
rect -3667 294349 -3549 294467
rect -3667 276509 -3549 276627
rect -3667 276349 -3549 276467
rect -3667 258509 -3549 258627
rect -3667 258349 -3549 258467
rect -3667 240509 -3549 240627
rect -3667 240349 -3549 240467
rect -3667 222509 -3549 222627
rect -3667 222349 -3549 222467
rect -3667 204509 -3549 204627
rect -3667 204349 -3549 204467
rect -3667 186509 -3549 186627
rect -3667 186349 -3549 186467
rect -3667 168509 -3549 168627
rect -3667 168349 -3549 168467
rect -3667 150509 -3549 150627
rect -3667 150349 -3549 150467
rect -3667 132509 -3549 132627
rect -3667 132349 -3549 132467
rect -3667 114509 -3549 114627
rect -3667 114349 -3549 114467
rect -3667 96509 -3549 96627
rect -3667 96349 -3549 96467
rect -3667 78509 -3549 78627
rect -3667 78349 -3549 78467
rect -3667 60509 -3549 60627
rect -3667 60349 -3549 60467
rect -3667 42509 -3549 42627
rect -3667 42349 -3549 42467
rect -3667 24509 -3549 24627
rect -3667 24349 -3549 24467
rect -3667 6509 -3549 6627
rect -3667 6349 -3549 6467
rect -3207 354601 -3089 354719
rect -3207 354441 -3089 354559
rect -3207 337709 -3089 337827
rect -3207 337549 -3089 337667
rect -3207 319709 -3089 319827
rect -3207 319549 -3089 319667
rect -3207 301709 -3089 301827
rect -3207 301549 -3089 301667
rect -3207 283709 -3089 283827
rect -3207 283549 -3089 283667
rect -3207 265709 -3089 265827
rect -3207 265549 -3089 265667
rect -3207 247709 -3089 247827
rect -3207 247549 -3089 247667
rect -3207 229709 -3089 229827
rect -3207 229549 -3089 229667
rect -3207 211709 -3089 211827
rect -3207 211549 -3089 211667
rect -3207 193709 -3089 193827
rect -3207 193549 -3089 193667
rect -3207 175709 -3089 175827
rect -3207 175549 -3089 175667
rect -3207 157709 -3089 157827
rect -3207 157549 -3089 157667
rect -3207 139709 -3089 139827
rect -3207 139549 -3089 139667
rect -3207 121709 -3089 121827
rect -3207 121549 -3089 121667
rect -3207 103709 -3089 103827
rect -3207 103549 -3089 103667
rect -3207 85709 -3089 85827
rect -3207 85549 -3089 85667
rect -3207 67709 -3089 67827
rect -3207 67549 -3089 67667
rect -3207 49709 -3089 49827
rect -3207 49549 -3089 49667
rect -3207 31709 -3089 31827
rect -3207 31549 -3089 31667
rect -3207 13709 -3089 13827
rect -3207 13549 -3089 13667
rect -2747 354141 -2629 354259
rect -2747 353981 -2629 354099
rect 4093 354141 4211 354259
rect 4093 353981 4211 354099
rect -2747 346709 -2629 346827
rect -2747 346549 -2629 346667
rect -2747 328709 -2629 328827
rect -2747 328549 -2629 328667
rect -2747 310709 -2629 310827
rect -2747 310549 -2629 310667
rect -2747 292709 -2629 292827
rect -2747 292549 -2629 292667
rect -2747 274709 -2629 274827
rect -2747 274549 -2629 274667
rect -2747 256709 -2629 256827
rect -2747 256549 -2629 256667
rect -2747 238709 -2629 238827
rect -2747 238549 -2629 238667
rect -2747 220709 -2629 220827
rect -2747 220549 -2629 220667
rect -2747 202709 -2629 202827
rect -2747 202549 -2629 202667
rect -2747 184709 -2629 184827
rect -2747 184549 -2629 184667
rect -2747 166709 -2629 166827
rect -2747 166549 -2629 166667
rect -2747 148709 -2629 148827
rect -2747 148549 -2629 148667
rect -2747 130709 -2629 130827
rect -2747 130549 -2629 130667
rect -2747 112709 -2629 112827
rect -2747 112549 -2629 112667
rect -2747 94709 -2629 94827
rect -2747 94549 -2629 94667
rect -2747 76709 -2629 76827
rect -2747 76549 -2629 76667
rect -2747 58709 -2629 58827
rect -2747 58549 -2629 58667
rect -2747 40709 -2629 40827
rect -2747 40549 -2629 40667
rect -2747 22709 -2629 22827
rect -2747 22549 -2629 22667
rect -2747 4709 -2629 4827
rect -2747 4549 -2629 4667
rect -2287 353681 -2169 353799
rect -2287 353521 -2169 353639
rect -2287 335909 -2169 336027
rect -2287 335749 -2169 335867
rect -2287 317909 -2169 318027
rect -2287 317749 -2169 317867
rect -2287 299909 -2169 300027
rect -2287 299749 -2169 299867
rect -2287 281909 -2169 282027
rect -2287 281749 -2169 281867
rect -2287 263909 -2169 264027
rect -2287 263749 -2169 263867
rect -2287 245909 -2169 246027
rect -2287 245749 -2169 245867
rect -2287 227909 -2169 228027
rect -2287 227749 -2169 227867
rect -2287 209909 -2169 210027
rect -2287 209749 -2169 209867
rect -2287 191909 -2169 192027
rect -2287 191749 -2169 191867
rect -2287 173909 -2169 174027
rect -2287 173749 -2169 173867
rect -2287 155909 -2169 156027
rect -2287 155749 -2169 155867
rect -2287 137909 -2169 138027
rect -2287 137749 -2169 137867
rect -2287 119909 -2169 120027
rect -2287 119749 -2169 119867
rect -2287 101909 -2169 102027
rect -2287 101749 -2169 101867
rect -2287 83909 -2169 84027
rect -2287 83749 -2169 83867
rect -2287 65909 -2169 66027
rect -2287 65749 -2169 65867
rect -2287 47909 -2169 48027
rect -2287 47749 -2169 47867
rect -2287 29909 -2169 30027
rect -2287 29749 -2169 29867
rect -2287 11909 -2169 12027
rect -2287 11749 -2169 11867
rect -1827 353221 -1709 353339
rect -1827 353061 -1709 353179
rect 2293 353221 2411 353339
rect 2293 353061 2411 353179
rect -1827 344909 -1709 345027
rect -1827 344749 -1709 344867
rect -1827 326909 -1709 327027
rect -1827 326749 -1709 326867
rect -1827 308909 -1709 309027
rect -1827 308749 -1709 308867
rect -1827 290909 -1709 291027
rect -1827 290749 -1709 290867
rect -1827 272909 -1709 273027
rect -1827 272749 -1709 272867
rect -1827 254909 -1709 255027
rect -1827 254749 -1709 254867
rect -1827 236909 -1709 237027
rect -1827 236749 -1709 236867
rect -1827 218909 -1709 219027
rect -1827 218749 -1709 218867
rect -1827 200909 -1709 201027
rect -1827 200749 -1709 200867
rect -1827 182909 -1709 183027
rect -1827 182749 -1709 182867
rect -1827 164909 -1709 165027
rect -1827 164749 -1709 164867
rect -1827 146909 -1709 147027
rect -1827 146749 -1709 146867
rect -1827 128909 -1709 129027
rect -1827 128749 -1709 128867
rect -1827 110909 -1709 111027
rect -1827 110749 -1709 110867
rect -1827 92909 -1709 93027
rect -1827 92749 -1709 92867
rect -1827 74909 -1709 75027
rect -1827 74749 -1709 74867
rect -1827 56909 -1709 57027
rect -1827 56749 -1709 56867
rect -1827 38909 -1709 39027
rect -1827 38749 -1709 38867
rect -1827 20909 -1709 21027
rect -1827 20749 -1709 20867
rect -1827 2909 -1709 3027
rect -1827 2749 -1709 2867
rect -1367 352761 -1249 352879
rect -1367 352601 -1249 352719
rect -1367 334109 -1249 334227
rect -1367 333949 -1249 334067
rect -1367 316109 -1249 316227
rect -1367 315949 -1249 316067
rect -1367 298109 -1249 298227
rect -1367 297949 -1249 298067
rect -1367 280109 -1249 280227
rect -1367 279949 -1249 280067
rect -1367 262109 -1249 262227
rect -1367 261949 -1249 262067
rect -1367 244109 -1249 244227
rect -1367 243949 -1249 244067
rect -1367 226109 -1249 226227
rect -1367 225949 -1249 226067
rect -1367 208109 -1249 208227
rect -1367 207949 -1249 208067
rect -1367 190109 -1249 190227
rect -1367 189949 -1249 190067
rect -1367 172109 -1249 172227
rect -1367 171949 -1249 172067
rect -1367 154109 -1249 154227
rect -1367 153949 -1249 154067
rect -1367 136109 -1249 136227
rect -1367 135949 -1249 136067
rect -1367 118109 -1249 118227
rect -1367 117949 -1249 118067
rect -1367 100109 -1249 100227
rect -1367 99949 -1249 100067
rect -1367 82109 -1249 82227
rect -1367 81949 -1249 82067
rect -1367 64109 -1249 64227
rect -1367 63949 -1249 64067
rect -1367 46109 -1249 46227
rect -1367 45949 -1249 46067
rect -1367 28109 -1249 28227
rect -1367 27949 -1249 28067
rect -1367 10109 -1249 10227
rect -1367 9949 -1249 10067
rect -907 352301 -789 352419
rect -907 352141 -789 352259
rect 493 352301 611 352419
rect 493 352141 611 352259
rect 14893 355521 15011 355639
rect 14893 355361 15011 355479
rect 13093 354601 13211 354719
rect 13093 354441 13211 354559
rect 11293 353681 11411 353799
rect 11293 353521 11411 353639
rect 9493 352761 9611 352879
rect 9493 352601 9611 352719
rect 23893 355061 24011 355179
rect 23893 354901 24011 355019
rect 22093 354141 22211 354259
rect 22093 353981 22211 354099
rect 20293 353221 20411 353339
rect 20293 353061 20411 353179
rect 18493 352301 18611 352419
rect 18493 352141 18611 352259
rect 32893 355521 33011 355639
rect 32893 355361 33011 355479
rect 31093 354601 31211 354719
rect 31093 354441 31211 354559
rect 29293 353681 29411 353799
rect 29293 353521 29411 353639
rect 27493 352761 27611 352879
rect 27493 352601 27611 352719
rect 41893 355061 42011 355179
rect 41893 354901 42011 355019
rect 40093 354141 40211 354259
rect 40093 353981 40211 354099
rect 38293 353221 38411 353339
rect 38293 353061 38411 353179
rect 36493 352301 36611 352419
rect 36493 352141 36611 352259
rect 50893 355521 51011 355639
rect 50893 355361 51011 355479
rect 49093 354601 49211 354719
rect 49093 354441 49211 354559
rect 47293 353681 47411 353799
rect 47293 353521 47411 353639
rect 45493 352761 45611 352879
rect 45493 352601 45611 352719
rect 59893 355061 60011 355179
rect 59893 354901 60011 355019
rect 58093 354141 58211 354259
rect 58093 353981 58211 354099
rect 56293 353221 56411 353339
rect 56293 353061 56411 353179
rect 54493 352301 54611 352419
rect 54493 352141 54611 352259
rect 68893 355521 69011 355639
rect 68893 355361 69011 355479
rect 67093 354601 67211 354719
rect 67093 354441 67211 354559
rect 65293 353681 65411 353799
rect 65293 353521 65411 353639
rect 63493 352761 63611 352879
rect 63493 352601 63611 352719
rect 77893 355061 78011 355179
rect 77893 354901 78011 355019
rect 76093 354141 76211 354259
rect 76093 353981 76211 354099
rect 74293 353221 74411 353339
rect 74293 353061 74411 353179
rect 72493 352301 72611 352419
rect 72493 352141 72611 352259
rect 86893 355521 87011 355639
rect 86893 355361 87011 355479
rect 85093 354601 85211 354719
rect 85093 354441 85211 354559
rect 83293 353681 83411 353799
rect 83293 353521 83411 353639
rect 81493 352761 81611 352879
rect 81493 352601 81611 352719
rect 95893 355061 96011 355179
rect 95893 354901 96011 355019
rect 94093 354141 94211 354259
rect 94093 353981 94211 354099
rect 92293 353221 92411 353339
rect 92293 353061 92411 353179
rect 90493 352301 90611 352419
rect 90493 352141 90611 352259
rect 104893 355521 105011 355639
rect 104893 355361 105011 355479
rect 103093 354601 103211 354719
rect 103093 354441 103211 354559
rect 101293 353681 101411 353799
rect 101293 353521 101411 353639
rect 99493 352761 99611 352879
rect 99493 352601 99611 352719
rect 113893 355061 114011 355179
rect 113893 354901 114011 355019
rect 112093 354141 112211 354259
rect 112093 353981 112211 354099
rect 110293 353221 110411 353339
rect 110293 353061 110411 353179
rect 108493 352301 108611 352419
rect 108493 352141 108611 352259
rect 122893 355521 123011 355639
rect 122893 355361 123011 355479
rect 121093 354601 121211 354719
rect 121093 354441 121211 354559
rect 119293 353681 119411 353799
rect 119293 353521 119411 353639
rect 117493 352761 117611 352879
rect 117493 352601 117611 352719
rect 131893 355061 132011 355179
rect 131893 354901 132011 355019
rect 130093 354141 130211 354259
rect 130093 353981 130211 354099
rect 128293 353221 128411 353339
rect 128293 353061 128411 353179
rect 126493 352301 126611 352419
rect 126493 352141 126611 352259
rect 140893 355521 141011 355639
rect 140893 355361 141011 355479
rect 139093 354601 139211 354719
rect 139093 354441 139211 354559
rect 137293 353681 137411 353799
rect 137293 353521 137411 353639
rect 135493 352761 135611 352879
rect 135493 352601 135611 352719
rect 149893 355061 150011 355179
rect 149893 354901 150011 355019
rect 148093 354141 148211 354259
rect 148093 353981 148211 354099
rect 146293 353221 146411 353339
rect 146293 353061 146411 353179
rect 144493 352301 144611 352419
rect 144493 352141 144611 352259
rect 158893 355521 159011 355639
rect 158893 355361 159011 355479
rect 157093 354601 157211 354719
rect 157093 354441 157211 354559
rect 155293 353681 155411 353799
rect 155293 353521 155411 353639
rect 153493 352761 153611 352879
rect 153493 352601 153611 352719
rect 167893 355061 168011 355179
rect 167893 354901 168011 355019
rect 166093 354141 166211 354259
rect 166093 353981 166211 354099
rect 164293 353221 164411 353339
rect 164293 353061 164411 353179
rect 162493 352301 162611 352419
rect 162493 352141 162611 352259
rect 176893 355521 177011 355639
rect 176893 355361 177011 355479
rect 175093 354601 175211 354719
rect 175093 354441 175211 354559
rect 173293 353681 173411 353799
rect 173293 353521 173411 353639
rect 171493 352761 171611 352879
rect 171493 352601 171611 352719
rect 185893 355061 186011 355179
rect 185893 354901 186011 355019
rect 184093 354141 184211 354259
rect 184093 353981 184211 354099
rect 182293 353221 182411 353339
rect 182293 353061 182411 353179
rect 180493 352301 180611 352419
rect 180493 352141 180611 352259
rect 194893 355521 195011 355639
rect 194893 355361 195011 355479
rect 193093 354601 193211 354719
rect 193093 354441 193211 354559
rect 191293 353681 191411 353799
rect 191293 353521 191411 353639
rect 189493 352761 189611 352879
rect 189493 352601 189611 352719
rect 203893 355061 204011 355179
rect 203893 354901 204011 355019
rect 202093 354141 202211 354259
rect 202093 353981 202211 354099
rect 200293 353221 200411 353339
rect 200293 353061 200411 353179
rect 198493 352301 198611 352419
rect 198493 352141 198611 352259
rect 212893 355521 213011 355639
rect 212893 355361 213011 355479
rect 211093 354601 211211 354719
rect 211093 354441 211211 354559
rect 209293 353681 209411 353799
rect 209293 353521 209411 353639
rect 207493 352761 207611 352879
rect 207493 352601 207611 352719
rect 221893 355061 222011 355179
rect 221893 354901 222011 355019
rect 220093 354141 220211 354259
rect 220093 353981 220211 354099
rect 218293 353221 218411 353339
rect 218293 353061 218411 353179
rect 216493 352301 216611 352419
rect 216493 352141 216611 352259
rect 230893 355521 231011 355639
rect 230893 355361 231011 355479
rect 229093 354601 229211 354719
rect 229093 354441 229211 354559
rect 227293 353681 227411 353799
rect 227293 353521 227411 353639
rect 225493 352761 225611 352879
rect 225493 352601 225611 352719
rect 239893 355061 240011 355179
rect 239893 354901 240011 355019
rect 238093 354141 238211 354259
rect 238093 353981 238211 354099
rect 236293 353221 236411 353339
rect 236293 353061 236411 353179
rect 234493 352301 234611 352419
rect 234493 352141 234611 352259
rect 248893 355521 249011 355639
rect 248893 355361 249011 355479
rect 247093 354601 247211 354719
rect 247093 354441 247211 354559
rect 245293 353681 245411 353799
rect 245293 353521 245411 353639
rect 243493 352761 243611 352879
rect 243493 352601 243611 352719
rect 257893 355061 258011 355179
rect 257893 354901 258011 355019
rect 256093 354141 256211 354259
rect 256093 353981 256211 354099
rect 254293 353221 254411 353339
rect 254293 353061 254411 353179
rect 252493 352301 252611 352419
rect 252493 352141 252611 352259
rect 266893 355521 267011 355639
rect 266893 355361 267011 355479
rect 265093 354601 265211 354719
rect 265093 354441 265211 354559
rect 263293 353681 263411 353799
rect 263293 353521 263411 353639
rect 261493 352761 261611 352879
rect 261493 352601 261611 352719
rect 275893 355061 276011 355179
rect 275893 354901 276011 355019
rect 274093 354141 274211 354259
rect 274093 353981 274211 354099
rect 272293 353221 272411 353339
rect 272293 353061 272411 353179
rect 270493 352301 270611 352419
rect 270493 352141 270611 352259
rect 284893 355521 285011 355639
rect 284893 355361 285011 355479
rect 283093 354601 283211 354719
rect 283093 354441 283211 354559
rect 281293 353681 281411 353799
rect 281293 353521 281411 353639
rect 279493 352761 279611 352879
rect 279493 352601 279611 352719
rect 295971 355521 296089 355639
rect 295971 355361 296089 355479
rect 295511 355061 295629 355179
rect 295511 354901 295629 355019
rect 295051 354601 295169 354719
rect 295051 354441 295169 354559
rect 294591 354141 294709 354259
rect 294591 353981 294709 354099
rect 294131 353681 294249 353799
rect 294131 353521 294249 353639
rect 290293 353221 290411 353339
rect 290293 353061 290411 353179
rect 288493 352301 288611 352419
rect 288493 352141 288611 352259
rect 293671 353221 293789 353339
rect 293671 353061 293789 353179
rect 293211 352761 293329 352879
rect 293211 352601 293329 352719
rect 292751 352301 292869 352419
rect 292751 352141 292869 352259
rect -907 343109 -789 343227
rect -907 342949 -789 343067
rect -907 325109 -789 325227
rect -907 324949 -789 325067
rect -907 307109 -789 307227
rect -907 306949 -789 307067
rect -907 289109 -789 289227
rect -907 288949 -789 289067
rect -907 271109 -789 271227
rect -907 270949 -789 271067
rect -907 253109 -789 253227
rect -907 252949 -789 253067
rect -907 235109 -789 235227
rect -907 234949 -789 235067
rect -907 217109 -789 217227
rect -907 216949 -789 217067
rect -907 199109 -789 199227
rect -907 198949 -789 199067
rect -907 181109 -789 181227
rect -907 180949 -789 181067
rect -907 163109 -789 163227
rect -907 162949 -789 163067
rect -907 145109 -789 145227
rect -907 144949 -789 145067
rect -907 127109 -789 127227
rect -907 126949 -789 127067
rect -907 109109 -789 109227
rect -907 108949 -789 109067
rect -907 91109 -789 91227
rect -907 90949 -789 91067
rect -907 73109 -789 73227
rect -907 72949 -789 73067
rect -907 55109 -789 55227
rect -907 54949 -789 55067
rect -907 37109 -789 37227
rect -907 36949 -789 37067
rect -907 19109 -789 19227
rect -907 18949 -789 19067
rect -907 1109 -789 1227
rect -907 949 -789 1067
rect 292751 343109 292869 343227
rect 292751 342949 292869 343067
rect 292751 325109 292869 325227
rect 292751 324949 292869 325067
rect 292751 307109 292869 307227
rect 292751 306949 292869 307067
rect 292751 289109 292869 289227
rect 292751 288949 292869 289067
rect 292751 271109 292869 271227
rect 292751 270949 292869 271067
rect 292751 253109 292869 253227
rect 292751 252949 292869 253067
rect 292751 235109 292869 235227
rect 292751 234949 292869 235067
rect 292751 217109 292869 217227
rect 292751 216949 292869 217067
rect 292751 199109 292869 199227
rect 292751 198949 292869 199067
rect 292751 181109 292869 181227
rect 292751 180949 292869 181067
rect 292751 163109 292869 163227
rect 292751 162949 292869 163067
rect 292751 145109 292869 145227
rect 292751 144949 292869 145067
rect 292751 127109 292869 127227
rect 292751 126949 292869 127067
rect 292751 109109 292869 109227
rect 292751 108949 292869 109067
rect 292751 91109 292869 91227
rect 292751 90949 292869 91067
rect 292751 73109 292869 73227
rect 292751 72949 292869 73067
rect 292751 55109 292869 55227
rect 292751 54949 292869 55067
rect 292751 37109 292869 37227
rect 292751 36949 292869 37067
rect 292751 19109 292869 19227
rect 292751 18949 292869 19067
rect 292751 1109 292869 1227
rect 292751 949 292869 1067
rect -907 -291 -789 -173
rect -907 -451 -789 -333
rect 493 -291 611 -173
rect 493 -451 611 -333
rect -1367 -751 -1249 -633
rect -1367 -911 -1249 -793
rect -1827 -1211 -1709 -1093
rect -1827 -1371 -1709 -1253
rect 2293 -1211 2411 -1093
rect 2293 -1371 2411 -1253
rect -2287 -1671 -2169 -1553
rect -2287 -1831 -2169 -1713
rect -2747 -2131 -2629 -2013
rect -2747 -2291 -2629 -2173
rect 4093 -2131 4211 -2013
rect 4093 -2291 4211 -2173
rect -3207 -2591 -3089 -2473
rect -3207 -2751 -3089 -2633
rect -3667 -3051 -3549 -2933
rect -3667 -3211 -3549 -3093
rect 9493 -751 9611 -633
rect 9493 -911 9611 -793
rect 11293 -1671 11411 -1553
rect 11293 -1831 11411 -1713
rect 13093 -2591 13211 -2473
rect 13093 -2751 13211 -2633
rect 5893 -3051 6011 -2933
rect 5893 -3211 6011 -3093
rect -4127 -3511 -4009 -3393
rect -4127 -3671 -4009 -3553
rect 18493 -291 18611 -173
rect 18493 -451 18611 -333
rect 20293 -1211 20411 -1093
rect 20293 -1371 20411 -1253
rect 22093 -2131 22211 -2013
rect 22093 -2291 22211 -2173
rect 14893 -3511 15011 -3393
rect 14893 -3671 15011 -3553
rect 27493 -751 27611 -633
rect 27493 -911 27611 -793
rect 29293 -1671 29411 -1553
rect 29293 -1831 29411 -1713
rect 31093 -2591 31211 -2473
rect 31093 -2751 31211 -2633
rect 23893 -3051 24011 -2933
rect 23893 -3211 24011 -3093
rect 36493 -291 36611 -173
rect 36493 -451 36611 -333
rect 38293 -1211 38411 -1093
rect 38293 -1371 38411 -1253
rect 40093 -2131 40211 -2013
rect 40093 -2291 40211 -2173
rect 32893 -3511 33011 -3393
rect 32893 -3671 33011 -3553
rect 45493 -751 45611 -633
rect 45493 -911 45611 -793
rect 47293 -1671 47411 -1553
rect 47293 -1831 47411 -1713
rect 49093 -2591 49211 -2473
rect 49093 -2751 49211 -2633
rect 41893 -3051 42011 -2933
rect 41893 -3211 42011 -3093
rect 54493 -291 54611 -173
rect 54493 -451 54611 -333
rect 56293 -1211 56411 -1093
rect 56293 -1371 56411 -1253
rect 58093 -2131 58211 -2013
rect 58093 -2291 58211 -2173
rect 50893 -3511 51011 -3393
rect 50893 -3671 51011 -3553
rect 63493 -751 63611 -633
rect 63493 -911 63611 -793
rect 65293 -1671 65411 -1553
rect 65293 -1831 65411 -1713
rect 67093 -2591 67211 -2473
rect 67093 -2751 67211 -2633
rect 59893 -3051 60011 -2933
rect 59893 -3211 60011 -3093
rect 72493 -291 72611 -173
rect 72493 -451 72611 -333
rect 74293 -1211 74411 -1093
rect 74293 -1371 74411 -1253
rect 76093 -2131 76211 -2013
rect 76093 -2291 76211 -2173
rect 68893 -3511 69011 -3393
rect 68893 -3671 69011 -3553
rect 81493 -751 81611 -633
rect 81493 -911 81611 -793
rect 83293 -1671 83411 -1553
rect 83293 -1831 83411 -1713
rect 85093 -2591 85211 -2473
rect 85093 -2751 85211 -2633
rect 77893 -3051 78011 -2933
rect 77893 -3211 78011 -3093
rect 90493 -291 90611 -173
rect 90493 -451 90611 -333
rect 92293 -1211 92411 -1093
rect 92293 -1371 92411 -1253
rect 94093 -2131 94211 -2013
rect 94093 -2291 94211 -2173
rect 86893 -3511 87011 -3393
rect 86893 -3671 87011 -3553
rect 99493 -751 99611 -633
rect 99493 -911 99611 -793
rect 101293 -1671 101411 -1553
rect 101293 -1831 101411 -1713
rect 103093 -2591 103211 -2473
rect 103093 -2751 103211 -2633
rect 95893 -3051 96011 -2933
rect 95893 -3211 96011 -3093
rect 108493 -291 108611 -173
rect 108493 -451 108611 -333
rect 110293 -1211 110411 -1093
rect 110293 -1371 110411 -1253
rect 112093 -2131 112211 -2013
rect 112093 -2291 112211 -2173
rect 104893 -3511 105011 -3393
rect 104893 -3671 105011 -3553
rect 117493 -751 117611 -633
rect 117493 -911 117611 -793
rect 119293 -1671 119411 -1553
rect 119293 -1831 119411 -1713
rect 121093 -2591 121211 -2473
rect 121093 -2751 121211 -2633
rect 113893 -3051 114011 -2933
rect 113893 -3211 114011 -3093
rect 126493 -291 126611 -173
rect 126493 -451 126611 -333
rect 128293 -1211 128411 -1093
rect 128293 -1371 128411 -1253
rect 130093 -2131 130211 -2013
rect 130093 -2291 130211 -2173
rect 122893 -3511 123011 -3393
rect 122893 -3671 123011 -3553
rect 135493 -751 135611 -633
rect 135493 -911 135611 -793
rect 137293 -1671 137411 -1553
rect 137293 -1831 137411 -1713
rect 139093 -2591 139211 -2473
rect 139093 -2751 139211 -2633
rect 131893 -3051 132011 -2933
rect 131893 -3211 132011 -3093
rect 144493 -291 144611 -173
rect 144493 -451 144611 -333
rect 146293 -1211 146411 -1093
rect 146293 -1371 146411 -1253
rect 148093 -2131 148211 -2013
rect 148093 -2291 148211 -2173
rect 140893 -3511 141011 -3393
rect 140893 -3671 141011 -3553
rect 153493 -751 153611 -633
rect 153493 -911 153611 -793
rect 155293 -1671 155411 -1553
rect 155293 -1831 155411 -1713
rect 157093 -2591 157211 -2473
rect 157093 -2751 157211 -2633
rect 149893 -3051 150011 -2933
rect 149893 -3211 150011 -3093
rect 162493 -291 162611 -173
rect 162493 -451 162611 -333
rect 164293 -1211 164411 -1093
rect 164293 -1371 164411 -1253
rect 166093 -2131 166211 -2013
rect 166093 -2291 166211 -2173
rect 158893 -3511 159011 -3393
rect 158893 -3671 159011 -3553
rect 171493 -751 171611 -633
rect 171493 -911 171611 -793
rect 173293 -1671 173411 -1553
rect 173293 -1831 173411 -1713
rect 175093 -2591 175211 -2473
rect 175093 -2751 175211 -2633
rect 167893 -3051 168011 -2933
rect 167893 -3211 168011 -3093
rect 180493 -291 180611 -173
rect 180493 -451 180611 -333
rect 182293 -1211 182411 -1093
rect 182293 -1371 182411 -1253
rect 184093 -2131 184211 -2013
rect 184093 -2291 184211 -2173
rect 176893 -3511 177011 -3393
rect 176893 -3671 177011 -3553
rect 189493 -751 189611 -633
rect 189493 -911 189611 -793
rect 191293 -1671 191411 -1553
rect 191293 -1831 191411 -1713
rect 193093 -2591 193211 -2473
rect 193093 -2751 193211 -2633
rect 185893 -3051 186011 -2933
rect 185893 -3211 186011 -3093
rect 198493 -291 198611 -173
rect 198493 -451 198611 -333
rect 200293 -1211 200411 -1093
rect 200293 -1371 200411 -1253
rect 202093 -2131 202211 -2013
rect 202093 -2291 202211 -2173
rect 194893 -3511 195011 -3393
rect 194893 -3671 195011 -3553
rect 207493 -751 207611 -633
rect 207493 -911 207611 -793
rect 209293 -1671 209411 -1553
rect 209293 -1831 209411 -1713
rect 211093 -2591 211211 -2473
rect 211093 -2751 211211 -2633
rect 203893 -3051 204011 -2933
rect 203893 -3211 204011 -3093
rect 216493 -291 216611 -173
rect 216493 -451 216611 -333
rect 218293 -1211 218411 -1093
rect 218293 -1371 218411 -1253
rect 220093 -2131 220211 -2013
rect 220093 -2291 220211 -2173
rect 212893 -3511 213011 -3393
rect 212893 -3671 213011 -3553
rect 225493 -751 225611 -633
rect 225493 -911 225611 -793
rect 227293 -1671 227411 -1553
rect 227293 -1831 227411 -1713
rect 229093 -2591 229211 -2473
rect 229093 -2751 229211 -2633
rect 221893 -3051 222011 -2933
rect 221893 -3211 222011 -3093
rect 234493 -291 234611 -173
rect 234493 -451 234611 -333
rect 236293 -1211 236411 -1093
rect 236293 -1371 236411 -1253
rect 238093 -2131 238211 -2013
rect 238093 -2291 238211 -2173
rect 230893 -3511 231011 -3393
rect 230893 -3671 231011 -3553
rect 243493 -751 243611 -633
rect 243493 -911 243611 -793
rect 245293 -1671 245411 -1553
rect 245293 -1831 245411 -1713
rect 247093 -2591 247211 -2473
rect 247093 -2751 247211 -2633
rect 239893 -3051 240011 -2933
rect 239893 -3211 240011 -3093
rect 252493 -291 252611 -173
rect 252493 -451 252611 -333
rect 254293 -1211 254411 -1093
rect 254293 -1371 254411 -1253
rect 256093 -2131 256211 -2013
rect 256093 -2291 256211 -2173
rect 248893 -3511 249011 -3393
rect 248893 -3671 249011 -3553
rect 261493 -751 261611 -633
rect 261493 -911 261611 -793
rect 263293 -1671 263411 -1553
rect 263293 -1831 263411 -1713
rect 265093 -2591 265211 -2473
rect 265093 -2751 265211 -2633
rect 257893 -3051 258011 -2933
rect 257893 -3211 258011 -3093
rect 270493 -291 270611 -173
rect 270493 -451 270611 -333
rect 272293 -1211 272411 -1093
rect 272293 -1371 272411 -1253
rect 274093 -2131 274211 -2013
rect 274093 -2291 274211 -2173
rect 266893 -3511 267011 -3393
rect 266893 -3671 267011 -3553
rect 279493 -751 279611 -633
rect 279493 -911 279611 -793
rect 281293 -1671 281411 -1553
rect 281293 -1831 281411 -1713
rect 283093 -2591 283211 -2473
rect 283093 -2751 283211 -2633
rect 275893 -3051 276011 -2933
rect 275893 -3211 276011 -3093
rect 288493 -291 288611 -173
rect 288493 -451 288611 -333
rect 292751 -291 292869 -173
rect 292751 -451 292869 -333
rect 293211 334109 293329 334227
rect 293211 333949 293329 334067
rect 293211 316109 293329 316227
rect 293211 315949 293329 316067
rect 293211 298109 293329 298227
rect 293211 297949 293329 298067
rect 293211 280109 293329 280227
rect 293211 279949 293329 280067
rect 293211 262109 293329 262227
rect 293211 261949 293329 262067
rect 293211 244109 293329 244227
rect 293211 243949 293329 244067
rect 293211 226109 293329 226227
rect 293211 225949 293329 226067
rect 293211 208109 293329 208227
rect 293211 207949 293329 208067
rect 293211 190109 293329 190227
rect 293211 189949 293329 190067
rect 293211 172109 293329 172227
rect 293211 171949 293329 172067
rect 293211 154109 293329 154227
rect 293211 153949 293329 154067
rect 293211 136109 293329 136227
rect 293211 135949 293329 136067
rect 293211 118109 293329 118227
rect 293211 117949 293329 118067
rect 293211 100109 293329 100227
rect 293211 99949 293329 100067
rect 293211 82109 293329 82227
rect 293211 81949 293329 82067
rect 293211 64109 293329 64227
rect 293211 63949 293329 64067
rect 293211 46109 293329 46227
rect 293211 45949 293329 46067
rect 293211 28109 293329 28227
rect 293211 27949 293329 28067
rect 293211 10109 293329 10227
rect 293211 9949 293329 10067
rect 293211 -751 293329 -633
rect 293211 -911 293329 -793
rect 293671 344909 293789 345027
rect 293671 344749 293789 344867
rect 293671 326909 293789 327027
rect 293671 326749 293789 326867
rect 293671 308909 293789 309027
rect 293671 308749 293789 308867
rect 293671 290909 293789 291027
rect 293671 290749 293789 290867
rect 293671 272909 293789 273027
rect 293671 272749 293789 272867
rect 293671 254909 293789 255027
rect 293671 254749 293789 254867
rect 293671 236909 293789 237027
rect 293671 236749 293789 236867
rect 293671 218909 293789 219027
rect 293671 218749 293789 218867
rect 293671 200909 293789 201027
rect 293671 200749 293789 200867
rect 293671 182909 293789 183027
rect 293671 182749 293789 182867
rect 293671 164909 293789 165027
rect 293671 164749 293789 164867
rect 293671 146909 293789 147027
rect 293671 146749 293789 146867
rect 293671 128909 293789 129027
rect 293671 128749 293789 128867
rect 293671 110909 293789 111027
rect 293671 110749 293789 110867
rect 293671 92909 293789 93027
rect 293671 92749 293789 92867
rect 293671 74909 293789 75027
rect 293671 74749 293789 74867
rect 293671 56909 293789 57027
rect 293671 56749 293789 56867
rect 293671 38909 293789 39027
rect 293671 38749 293789 38867
rect 293671 20909 293789 21027
rect 293671 20749 293789 20867
rect 293671 2909 293789 3027
rect 293671 2749 293789 2867
rect 290293 -1211 290411 -1093
rect 290293 -1371 290411 -1253
rect 293671 -1211 293789 -1093
rect 293671 -1371 293789 -1253
rect 294131 335909 294249 336027
rect 294131 335749 294249 335867
rect 294131 317909 294249 318027
rect 294131 317749 294249 317867
rect 294131 299909 294249 300027
rect 294131 299749 294249 299867
rect 294131 281909 294249 282027
rect 294131 281749 294249 281867
rect 294131 263909 294249 264027
rect 294131 263749 294249 263867
rect 294131 245909 294249 246027
rect 294131 245749 294249 245867
rect 294131 227909 294249 228027
rect 294131 227749 294249 227867
rect 294131 209909 294249 210027
rect 294131 209749 294249 209867
rect 294131 191909 294249 192027
rect 294131 191749 294249 191867
rect 294131 173909 294249 174027
rect 294131 173749 294249 173867
rect 294131 155909 294249 156027
rect 294131 155749 294249 155867
rect 294131 137909 294249 138027
rect 294131 137749 294249 137867
rect 294131 119909 294249 120027
rect 294131 119749 294249 119867
rect 294131 101909 294249 102027
rect 294131 101749 294249 101867
rect 294131 83909 294249 84027
rect 294131 83749 294249 83867
rect 294131 65909 294249 66027
rect 294131 65749 294249 65867
rect 294131 47909 294249 48027
rect 294131 47749 294249 47867
rect 294131 29909 294249 30027
rect 294131 29749 294249 29867
rect 294131 11909 294249 12027
rect 294131 11749 294249 11867
rect 294131 -1671 294249 -1553
rect 294131 -1831 294249 -1713
rect 294591 346709 294709 346827
rect 294591 346549 294709 346667
rect 294591 328709 294709 328827
rect 294591 328549 294709 328667
rect 294591 310709 294709 310827
rect 294591 310549 294709 310667
rect 294591 292709 294709 292827
rect 294591 292549 294709 292667
rect 294591 274709 294709 274827
rect 294591 274549 294709 274667
rect 294591 256709 294709 256827
rect 294591 256549 294709 256667
rect 294591 238709 294709 238827
rect 294591 238549 294709 238667
rect 294591 220709 294709 220827
rect 294591 220549 294709 220667
rect 294591 202709 294709 202827
rect 294591 202549 294709 202667
rect 294591 184709 294709 184827
rect 294591 184549 294709 184667
rect 294591 166709 294709 166827
rect 294591 166549 294709 166667
rect 294591 148709 294709 148827
rect 294591 148549 294709 148667
rect 294591 130709 294709 130827
rect 294591 130549 294709 130667
rect 294591 112709 294709 112827
rect 294591 112549 294709 112667
rect 294591 94709 294709 94827
rect 294591 94549 294709 94667
rect 294591 76709 294709 76827
rect 294591 76549 294709 76667
rect 294591 58709 294709 58827
rect 294591 58549 294709 58667
rect 294591 40709 294709 40827
rect 294591 40549 294709 40667
rect 294591 22709 294709 22827
rect 294591 22549 294709 22667
rect 294591 4709 294709 4827
rect 294591 4549 294709 4667
rect 294591 -2131 294709 -2013
rect 294591 -2291 294709 -2173
rect 295051 337709 295169 337827
rect 295051 337549 295169 337667
rect 295051 319709 295169 319827
rect 295051 319549 295169 319667
rect 295051 301709 295169 301827
rect 295051 301549 295169 301667
rect 295051 283709 295169 283827
rect 295051 283549 295169 283667
rect 295051 265709 295169 265827
rect 295051 265549 295169 265667
rect 295051 247709 295169 247827
rect 295051 247549 295169 247667
rect 295051 229709 295169 229827
rect 295051 229549 295169 229667
rect 295051 211709 295169 211827
rect 295051 211549 295169 211667
rect 295051 193709 295169 193827
rect 295051 193549 295169 193667
rect 295051 175709 295169 175827
rect 295051 175549 295169 175667
rect 295051 157709 295169 157827
rect 295051 157549 295169 157667
rect 295051 139709 295169 139827
rect 295051 139549 295169 139667
rect 295051 121709 295169 121827
rect 295051 121549 295169 121667
rect 295051 103709 295169 103827
rect 295051 103549 295169 103667
rect 295051 85709 295169 85827
rect 295051 85549 295169 85667
rect 295051 67709 295169 67827
rect 295051 67549 295169 67667
rect 295051 49709 295169 49827
rect 295051 49549 295169 49667
rect 295051 31709 295169 31827
rect 295051 31549 295169 31667
rect 295051 13709 295169 13827
rect 295051 13549 295169 13667
rect 295051 -2591 295169 -2473
rect 295051 -2751 295169 -2633
rect 295511 348509 295629 348627
rect 295511 348349 295629 348467
rect 295511 330509 295629 330627
rect 295511 330349 295629 330467
rect 295511 312509 295629 312627
rect 295511 312349 295629 312467
rect 295511 294509 295629 294627
rect 295511 294349 295629 294467
rect 295511 276509 295629 276627
rect 295511 276349 295629 276467
rect 295511 258509 295629 258627
rect 295511 258349 295629 258467
rect 295511 240509 295629 240627
rect 295511 240349 295629 240467
rect 295511 222509 295629 222627
rect 295511 222349 295629 222467
rect 295511 204509 295629 204627
rect 295511 204349 295629 204467
rect 295511 186509 295629 186627
rect 295511 186349 295629 186467
rect 295511 168509 295629 168627
rect 295511 168349 295629 168467
rect 295511 150509 295629 150627
rect 295511 150349 295629 150467
rect 295511 132509 295629 132627
rect 295511 132349 295629 132467
rect 295511 114509 295629 114627
rect 295511 114349 295629 114467
rect 295511 96509 295629 96627
rect 295511 96349 295629 96467
rect 295511 78509 295629 78627
rect 295511 78349 295629 78467
rect 295511 60509 295629 60627
rect 295511 60349 295629 60467
rect 295511 42509 295629 42627
rect 295511 42349 295629 42467
rect 295511 24509 295629 24627
rect 295511 24349 295629 24467
rect 295511 6509 295629 6627
rect 295511 6349 295629 6467
rect 295511 -3051 295629 -2933
rect 295511 -3211 295629 -3093
rect 295971 339509 296089 339627
rect 295971 339349 296089 339467
rect 295971 321509 296089 321627
rect 295971 321349 296089 321467
rect 295971 303509 296089 303627
rect 295971 303349 296089 303467
rect 295971 285509 296089 285627
rect 295971 285349 296089 285467
rect 295971 267509 296089 267627
rect 295971 267349 296089 267467
rect 295971 249509 296089 249627
rect 295971 249349 296089 249467
rect 295971 231509 296089 231627
rect 295971 231349 296089 231467
rect 295971 213509 296089 213627
rect 295971 213349 296089 213467
rect 295971 195509 296089 195627
rect 295971 195349 296089 195467
rect 295971 177509 296089 177627
rect 295971 177349 296089 177467
rect 295971 159509 296089 159627
rect 295971 159349 296089 159467
rect 295971 141509 296089 141627
rect 295971 141349 296089 141467
rect 295971 123509 296089 123627
rect 295971 123349 296089 123467
rect 295971 105509 296089 105627
rect 295971 105349 296089 105467
rect 295971 87509 296089 87627
rect 295971 87349 296089 87467
rect 295971 69509 296089 69627
rect 295971 69349 296089 69467
rect 295971 51509 296089 51627
rect 295971 51349 296089 51467
rect 295971 33509 296089 33627
rect 295971 33349 296089 33467
rect 295971 15509 296089 15627
rect 295971 15349 296089 15467
rect 284893 -3511 285011 -3393
rect 284893 -3671 285011 -3553
rect 295971 -3511 296089 -3393
rect 295971 -3671 296089 -3553
<< metal5 >>
rect -4218 355650 -3918 355651
rect 14802 355650 15102 355651
rect 32802 355650 33102 355651
rect 50802 355650 51102 355651
rect 68802 355650 69102 355651
rect 86802 355650 87102 355651
rect 104802 355650 105102 355651
rect 122802 355650 123102 355651
rect 140802 355650 141102 355651
rect 158802 355650 159102 355651
rect 176802 355650 177102 355651
rect 194802 355650 195102 355651
rect 212802 355650 213102 355651
rect 230802 355650 231102 355651
rect 248802 355650 249102 355651
rect 266802 355650 267102 355651
rect 284802 355650 285102 355651
rect 295880 355650 296180 355651
rect -4218 355639 296180 355650
rect -4218 355521 -4127 355639
rect -4009 355521 14893 355639
rect 15011 355521 32893 355639
rect 33011 355521 50893 355639
rect 51011 355521 68893 355639
rect 69011 355521 86893 355639
rect 87011 355521 104893 355639
rect 105011 355521 122893 355639
rect 123011 355521 140893 355639
rect 141011 355521 158893 355639
rect 159011 355521 176893 355639
rect 177011 355521 194893 355639
rect 195011 355521 212893 355639
rect 213011 355521 230893 355639
rect 231011 355521 248893 355639
rect 249011 355521 266893 355639
rect 267011 355521 284893 355639
rect 285011 355521 295971 355639
rect 296089 355521 296180 355639
rect -4218 355479 296180 355521
rect -4218 355361 -4127 355479
rect -4009 355361 14893 355479
rect 15011 355361 32893 355479
rect 33011 355361 50893 355479
rect 51011 355361 68893 355479
rect 69011 355361 86893 355479
rect 87011 355361 104893 355479
rect 105011 355361 122893 355479
rect 123011 355361 140893 355479
rect 141011 355361 158893 355479
rect 159011 355361 176893 355479
rect 177011 355361 194893 355479
rect 195011 355361 212893 355479
rect 213011 355361 230893 355479
rect 231011 355361 248893 355479
rect 249011 355361 266893 355479
rect 267011 355361 284893 355479
rect 285011 355361 295971 355479
rect 296089 355361 296180 355479
rect -4218 355350 296180 355361
rect -4218 355349 -3918 355350
rect 14802 355349 15102 355350
rect 32802 355349 33102 355350
rect 50802 355349 51102 355350
rect 68802 355349 69102 355350
rect 86802 355349 87102 355350
rect 104802 355349 105102 355350
rect 122802 355349 123102 355350
rect 140802 355349 141102 355350
rect 158802 355349 159102 355350
rect 176802 355349 177102 355350
rect 194802 355349 195102 355350
rect 212802 355349 213102 355350
rect 230802 355349 231102 355350
rect 248802 355349 249102 355350
rect 266802 355349 267102 355350
rect 284802 355349 285102 355350
rect 295880 355349 296180 355350
rect -3758 355190 -3458 355191
rect 5802 355190 6102 355191
rect 23802 355190 24102 355191
rect 41802 355190 42102 355191
rect 59802 355190 60102 355191
rect 77802 355190 78102 355191
rect 95802 355190 96102 355191
rect 113802 355190 114102 355191
rect 131802 355190 132102 355191
rect 149802 355190 150102 355191
rect 167802 355190 168102 355191
rect 185802 355190 186102 355191
rect 203802 355190 204102 355191
rect 221802 355190 222102 355191
rect 239802 355190 240102 355191
rect 257802 355190 258102 355191
rect 275802 355190 276102 355191
rect 295420 355190 295720 355191
rect -3758 355179 295720 355190
rect -3758 355061 -3667 355179
rect -3549 355061 5893 355179
rect 6011 355061 23893 355179
rect 24011 355061 41893 355179
rect 42011 355061 59893 355179
rect 60011 355061 77893 355179
rect 78011 355061 95893 355179
rect 96011 355061 113893 355179
rect 114011 355061 131893 355179
rect 132011 355061 149893 355179
rect 150011 355061 167893 355179
rect 168011 355061 185893 355179
rect 186011 355061 203893 355179
rect 204011 355061 221893 355179
rect 222011 355061 239893 355179
rect 240011 355061 257893 355179
rect 258011 355061 275893 355179
rect 276011 355061 295511 355179
rect 295629 355061 295720 355179
rect -3758 355019 295720 355061
rect -3758 354901 -3667 355019
rect -3549 354901 5893 355019
rect 6011 354901 23893 355019
rect 24011 354901 41893 355019
rect 42011 354901 59893 355019
rect 60011 354901 77893 355019
rect 78011 354901 95893 355019
rect 96011 354901 113893 355019
rect 114011 354901 131893 355019
rect 132011 354901 149893 355019
rect 150011 354901 167893 355019
rect 168011 354901 185893 355019
rect 186011 354901 203893 355019
rect 204011 354901 221893 355019
rect 222011 354901 239893 355019
rect 240011 354901 257893 355019
rect 258011 354901 275893 355019
rect 276011 354901 295511 355019
rect 295629 354901 295720 355019
rect -3758 354890 295720 354901
rect -3758 354889 -3458 354890
rect 5802 354889 6102 354890
rect 23802 354889 24102 354890
rect 41802 354889 42102 354890
rect 59802 354889 60102 354890
rect 77802 354889 78102 354890
rect 95802 354889 96102 354890
rect 113802 354889 114102 354890
rect 131802 354889 132102 354890
rect 149802 354889 150102 354890
rect 167802 354889 168102 354890
rect 185802 354889 186102 354890
rect 203802 354889 204102 354890
rect 221802 354889 222102 354890
rect 239802 354889 240102 354890
rect 257802 354889 258102 354890
rect 275802 354889 276102 354890
rect 295420 354889 295720 354890
rect -3298 354730 -2998 354731
rect 13002 354730 13302 354731
rect 31002 354730 31302 354731
rect 49002 354730 49302 354731
rect 67002 354730 67302 354731
rect 85002 354730 85302 354731
rect 103002 354730 103302 354731
rect 121002 354730 121302 354731
rect 139002 354730 139302 354731
rect 157002 354730 157302 354731
rect 175002 354730 175302 354731
rect 193002 354730 193302 354731
rect 211002 354730 211302 354731
rect 229002 354730 229302 354731
rect 247002 354730 247302 354731
rect 265002 354730 265302 354731
rect 283002 354730 283302 354731
rect 294960 354730 295260 354731
rect -3298 354719 295260 354730
rect -3298 354601 -3207 354719
rect -3089 354601 13093 354719
rect 13211 354601 31093 354719
rect 31211 354601 49093 354719
rect 49211 354601 67093 354719
rect 67211 354601 85093 354719
rect 85211 354601 103093 354719
rect 103211 354601 121093 354719
rect 121211 354601 139093 354719
rect 139211 354601 157093 354719
rect 157211 354601 175093 354719
rect 175211 354601 193093 354719
rect 193211 354601 211093 354719
rect 211211 354601 229093 354719
rect 229211 354601 247093 354719
rect 247211 354601 265093 354719
rect 265211 354601 283093 354719
rect 283211 354601 295051 354719
rect 295169 354601 295260 354719
rect -3298 354559 295260 354601
rect -3298 354441 -3207 354559
rect -3089 354441 13093 354559
rect 13211 354441 31093 354559
rect 31211 354441 49093 354559
rect 49211 354441 67093 354559
rect 67211 354441 85093 354559
rect 85211 354441 103093 354559
rect 103211 354441 121093 354559
rect 121211 354441 139093 354559
rect 139211 354441 157093 354559
rect 157211 354441 175093 354559
rect 175211 354441 193093 354559
rect 193211 354441 211093 354559
rect 211211 354441 229093 354559
rect 229211 354441 247093 354559
rect 247211 354441 265093 354559
rect 265211 354441 283093 354559
rect 283211 354441 295051 354559
rect 295169 354441 295260 354559
rect -3298 354430 295260 354441
rect -3298 354429 -2998 354430
rect 13002 354429 13302 354430
rect 31002 354429 31302 354430
rect 49002 354429 49302 354430
rect 67002 354429 67302 354430
rect 85002 354429 85302 354430
rect 103002 354429 103302 354430
rect 121002 354429 121302 354430
rect 139002 354429 139302 354430
rect 157002 354429 157302 354430
rect 175002 354429 175302 354430
rect 193002 354429 193302 354430
rect 211002 354429 211302 354430
rect 229002 354429 229302 354430
rect 247002 354429 247302 354430
rect 265002 354429 265302 354430
rect 283002 354429 283302 354430
rect 294960 354429 295260 354430
rect -2838 354270 -2538 354271
rect 4002 354270 4302 354271
rect 22002 354270 22302 354271
rect 40002 354270 40302 354271
rect 58002 354270 58302 354271
rect 76002 354270 76302 354271
rect 94002 354270 94302 354271
rect 112002 354270 112302 354271
rect 130002 354270 130302 354271
rect 148002 354270 148302 354271
rect 166002 354270 166302 354271
rect 184002 354270 184302 354271
rect 202002 354270 202302 354271
rect 220002 354270 220302 354271
rect 238002 354270 238302 354271
rect 256002 354270 256302 354271
rect 274002 354270 274302 354271
rect 294500 354270 294800 354271
rect -2838 354259 294800 354270
rect -2838 354141 -2747 354259
rect -2629 354141 4093 354259
rect 4211 354141 22093 354259
rect 22211 354141 40093 354259
rect 40211 354141 58093 354259
rect 58211 354141 76093 354259
rect 76211 354141 94093 354259
rect 94211 354141 112093 354259
rect 112211 354141 130093 354259
rect 130211 354141 148093 354259
rect 148211 354141 166093 354259
rect 166211 354141 184093 354259
rect 184211 354141 202093 354259
rect 202211 354141 220093 354259
rect 220211 354141 238093 354259
rect 238211 354141 256093 354259
rect 256211 354141 274093 354259
rect 274211 354141 294591 354259
rect 294709 354141 294800 354259
rect -2838 354099 294800 354141
rect -2838 353981 -2747 354099
rect -2629 353981 4093 354099
rect 4211 353981 22093 354099
rect 22211 353981 40093 354099
rect 40211 353981 58093 354099
rect 58211 353981 76093 354099
rect 76211 353981 94093 354099
rect 94211 353981 112093 354099
rect 112211 353981 130093 354099
rect 130211 353981 148093 354099
rect 148211 353981 166093 354099
rect 166211 353981 184093 354099
rect 184211 353981 202093 354099
rect 202211 353981 220093 354099
rect 220211 353981 238093 354099
rect 238211 353981 256093 354099
rect 256211 353981 274093 354099
rect 274211 353981 294591 354099
rect 294709 353981 294800 354099
rect -2838 353970 294800 353981
rect -2838 353969 -2538 353970
rect 4002 353969 4302 353970
rect 22002 353969 22302 353970
rect 40002 353969 40302 353970
rect 58002 353969 58302 353970
rect 76002 353969 76302 353970
rect 94002 353969 94302 353970
rect 112002 353969 112302 353970
rect 130002 353969 130302 353970
rect 148002 353969 148302 353970
rect 166002 353969 166302 353970
rect 184002 353969 184302 353970
rect 202002 353969 202302 353970
rect 220002 353969 220302 353970
rect 238002 353969 238302 353970
rect 256002 353969 256302 353970
rect 274002 353969 274302 353970
rect 294500 353969 294800 353970
rect -2378 353810 -2078 353811
rect 11202 353810 11502 353811
rect 29202 353810 29502 353811
rect 47202 353810 47502 353811
rect 65202 353810 65502 353811
rect 83202 353810 83502 353811
rect 101202 353810 101502 353811
rect 119202 353810 119502 353811
rect 137202 353810 137502 353811
rect 155202 353810 155502 353811
rect 173202 353810 173502 353811
rect 191202 353810 191502 353811
rect 209202 353810 209502 353811
rect 227202 353810 227502 353811
rect 245202 353810 245502 353811
rect 263202 353810 263502 353811
rect 281202 353810 281502 353811
rect 294040 353810 294340 353811
rect -2378 353799 294340 353810
rect -2378 353681 -2287 353799
rect -2169 353681 11293 353799
rect 11411 353681 29293 353799
rect 29411 353681 47293 353799
rect 47411 353681 65293 353799
rect 65411 353681 83293 353799
rect 83411 353681 101293 353799
rect 101411 353681 119293 353799
rect 119411 353681 137293 353799
rect 137411 353681 155293 353799
rect 155411 353681 173293 353799
rect 173411 353681 191293 353799
rect 191411 353681 209293 353799
rect 209411 353681 227293 353799
rect 227411 353681 245293 353799
rect 245411 353681 263293 353799
rect 263411 353681 281293 353799
rect 281411 353681 294131 353799
rect 294249 353681 294340 353799
rect -2378 353639 294340 353681
rect -2378 353521 -2287 353639
rect -2169 353521 11293 353639
rect 11411 353521 29293 353639
rect 29411 353521 47293 353639
rect 47411 353521 65293 353639
rect 65411 353521 83293 353639
rect 83411 353521 101293 353639
rect 101411 353521 119293 353639
rect 119411 353521 137293 353639
rect 137411 353521 155293 353639
rect 155411 353521 173293 353639
rect 173411 353521 191293 353639
rect 191411 353521 209293 353639
rect 209411 353521 227293 353639
rect 227411 353521 245293 353639
rect 245411 353521 263293 353639
rect 263411 353521 281293 353639
rect 281411 353521 294131 353639
rect 294249 353521 294340 353639
rect -2378 353510 294340 353521
rect -2378 353509 -2078 353510
rect 11202 353509 11502 353510
rect 29202 353509 29502 353510
rect 47202 353509 47502 353510
rect 65202 353509 65502 353510
rect 83202 353509 83502 353510
rect 101202 353509 101502 353510
rect 119202 353509 119502 353510
rect 137202 353509 137502 353510
rect 155202 353509 155502 353510
rect 173202 353509 173502 353510
rect 191202 353509 191502 353510
rect 209202 353509 209502 353510
rect 227202 353509 227502 353510
rect 245202 353509 245502 353510
rect 263202 353509 263502 353510
rect 281202 353509 281502 353510
rect 294040 353509 294340 353510
rect -1918 353350 -1618 353351
rect 2202 353350 2502 353351
rect 20202 353350 20502 353351
rect 38202 353350 38502 353351
rect 56202 353350 56502 353351
rect 74202 353350 74502 353351
rect 92202 353350 92502 353351
rect 110202 353350 110502 353351
rect 128202 353350 128502 353351
rect 146202 353350 146502 353351
rect 164202 353350 164502 353351
rect 182202 353350 182502 353351
rect 200202 353350 200502 353351
rect 218202 353350 218502 353351
rect 236202 353350 236502 353351
rect 254202 353350 254502 353351
rect 272202 353350 272502 353351
rect 290202 353350 290502 353351
rect 293580 353350 293880 353351
rect -1918 353339 293880 353350
rect -1918 353221 -1827 353339
rect -1709 353221 2293 353339
rect 2411 353221 20293 353339
rect 20411 353221 38293 353339
rect 38411 353221 56293 353339
rect 56411 353221 74293 353339
rect 74411 353221 92293 353339
rect 92411 353221 110293 353339
rect 110411 353221 128293 353339
rect 128411 353221 146293 353339
rect 146411 353221 164293 353339
rect 164411 353221 182293 353339
rect 182411 353221 200293 353339
rect 200411 353221 218293 353339
rect 218411 353221 236293 353339
rect 236411 353221 254293 353339
rect 254411 353221 272293 353339
rect 272411 353221 290293 353339
rect 290411 353221 293671 353339
rect 293789 353221 293880 353339
rect -1918 353179 293880 353221
rect -1918 353061 -1827 353179
rect -1709 353061 2293 353179
rect 2411 353061 20293 353179
rect 20411 353061 38293 353179
rect 38411 353061 56293 353179
rect 56411 353061 74293 353179
rect 74411 353061 92293 353179
rect 92411 353061 110293 353179
rect 110411 353061 128293 353179
rect 128411 353061 146293 353179
rect 146411 353061 164293 353179
rect 164411 353061 182293 353179
rect 182411 353061 200293 353179
rect 200411 353061 218293 353179
rect 218411 353061 236293 353179
rect 236411 353061 254293 353179
rect 254411 353061 272293 353179
rect 272411 353061 290293 353179
rect 290411 353061 293671 353179
rect 293789 353061 293880 353179
rect -1918 353050 293880 353061
rect -1918 353049 -1618 353050
rect 2202 353049 2502 353050
rect 20202 353049 20502 353050
rect 38202 353049 38502 353050
rect 56202 353049 56502 353050
rect 74202 353049 74502 353050
rect 92202 353049 92502 353050
rect 110202 353049 110502 353050
rect 128202 353049 128502 353050
rect 146202 353049 146502 353050
rect 164202 353049 164502 353050
rect 182202 353049 182502 353050
rect 200202 353049 200502 353050
rect 218202 353049 218502 353050
rect 236202 353049 236502 353050
rect 254202 353049 254502 353050
rect 272202 353049 272502 353050
rect 290202 353049 290502 353050
rect 293580 353049 293880 353050
rect -1458 352890 -1158 352891
rect 9402 352890 9702 352891
rect 27402 352890 27702 352891
rect 45402 352890 45702 352891
rect 63402 352890 63702 352891
rect 81402 352890 81702 352891
rect 99402 352890 99702 352891
rect 117402 352890 117702 352891
rect 135402 352890 135702 352891
rect 153402 352890 153702 352891
rect 171402 352890 171702 352891
rect 189402 352890 189702 352891
rect 207402 352890 207702 352891
rect 225402 352890 225702 352891
rect 243402 352890 243702 352891
rect 261402 352890 261702 352891
rect 279402 352890 279702 352891
rect 293120 352890 293420 352891
rect -1458 352879 293420 352890
rect -1458 352761 -1367 352879
rect -1249 352761 9493 352879
rect 9611 352761 27493 352879
rect 27611 352761 45493 352879
rect 45611 352761 63493 352879
rect 63611 352761 81493 352879
rect 81611 352761 99493 352879
rect 99611 352761 117493 352879
rect 117611 352761 135493 352879
rect 135611 352761 153493 352879
rect 153611 352761 171493 352879
rect 171611 352761 189493 352879
rect 189611 352761 207493 352879
rect 207611 352761 225493 352879
rect 225611 352761 243493 352879
rect 243611 352761 261493 352879
rect 261611 352761 279493 352879
rect 279611 352761 293211 352879
rect 293329 352761 293420 352879
rect -1458 352719 293420 352761
rect -1458 352601 -1367 352719
rect -1249 352601 9493 352719
rect 9611 352601 27493 352719
rect 27611 352601 45493 352719
rect 45611 352601 63493 352719
rect 63611 352601 81493 352719
rect 81611 352601 99493 352719
rect 99611 352601 117493 352719
rect 117611 352601 135493 352719
rect 135611 352601 153493 352719
rect 153611 352601 171493 352719
rect 171611 352601 189493 352719
rect 189611 352601 207493 352719
rect 207611 352601 225493 352719
rect 225611 352601 243493 352719
rect 243611 352601 261493 352719
rect 261611 352601 279493 352719
rect 279611 352601 293211 352719
rect 293329 352601 293420 352719
rect -1458 352590 293420 352601
rect -1458 352589 -1158 352590
rect 9402 352589 9702 352590
rect 27402 352589 27702 352590
rect 45402 352589 45702 352590
rect 63402 352589 63702 352590
rect 81402 352589 81702 352590
rect 99402 352589 99702 352590
rect 117402 352589 117702 352590
rect 135402 352589 135702 352590
rect 153402 352589 153702 352590
rect 171402 352589 171702 352590
rect 189402 352589 189702 352590
rect 207402 352589 207702 352590
rect 225402 352589 225702 352590
rect 243402 352589 243702 352590
rect 261402 352589 261702 352590
rect 279402 352589 279702 352590
rect 293120 352589 293420 352590
rect -998 352430 -698 352431
rect 402 352430 702 352431
rect 18402 352430 18702 352431
rect 36402 352430 36702 352431
rect 54402 352430 54702 352431
rect 72402 352430 72702 352431
rect 90402 352430 90702 352431
rect 108402 352430 108702 352431
rect 126402 352430 126702 352431
rect 144402 352430 144702 352431
rect 162402 352430 162702 352431
rect 180402 352430 180702 352431
rect 198402 352430 198702 352431
rect 216402 352430 216702 352431
rect 234402 352430 234702 352431
rect 252402 352430 252702 352431
rect 270402 352430 270702 352431
rect 288402 352430 288702 352431
rect 292660 352430 292960 352431
rect -998 352419 292960 352430
rect -998 352301 -907 352419
rect -789 352301 493 352419
rect 611 352301 18493 352419
rect 18611 352301 36493 352419
rect 36611 352301 54493 352419
rect 54611 352301 72493 352419
rect 72611 352301 90493 352419
rect 90611 352301 108493 352419
rect 108611 352301 126493 352419
rect 126611 352301 144493 352419
rect 144611 352301 162493 352419
rect 162611 352301 180493 352419
rect 180611 352301 198493 352419
rect 198611 352301 216493 352419
rect 216611 352301 234493 352419
rect 234611 352301 252493 352419
rect 252611 352301 270493 352419
rect 270611 352301 288493 352419
rect 288611 352301 292751 352419
rect 292869 352301 292960 352419
rect -998 352259 292960 352301
rect -998 352141 -907 352259
rect -789 352141 493 352259
rect 611 352141 18493 352259
rect 18611 352141 36493 352259
rect 36611 352141 54493 352259
rect 54611 352141 72493 352259
rect 72611 352141 90493 352259
rect 90611 352141 108493 352259
rect 108611 352141 126493 352259
rect 126611 352141 144493 352259
rect 144611 352141 162493 352259
rect 162611 352141 180493 352259
rect 180611 352141 198493 352259
rect 198611 352141 216493 352259
rect 216611 352141 234493 352259
rect 234611 352141 252493 352259
rect 252611 352141 270493 352259
rect 270611 352141 288493 352259
rect 288611 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 352130 292960 352141
rect -998 352129 -698 352130
rect 402 352129 702 352130
rect 18402 352129 18702 352130
rect 36402 352129 36702 352130
rect 54402 352129 54702 352130
rect 72402 352129 72702 352130
rect 90402 352129 90702 352130
rect 108402 352129 108702 352130
rect 126402 352129 126702 352130
rect 144402 352129 144702 352130
rect 162402 352129 162702 352130
rect 180402 352129 180702 352130
rect 198402 352129 198702 352130
rect 216402 352129 216702 352130
rect 234402 352129 234702 352130
rect 252402 352129 252702 352130
rect 270402 352129 270702 352130
rect 288402 352129 288702 352130
rect 292660 352129 292960 352130
rect -3758 348638 -3458 348639
rect 295420 348638 295720 348639
rect -4218 348627 240 348638
rect -4218 348509 -3667 348627
rect -3549 348509 240 348627
rect -4218 348467 240 348509
rect -4218 348349 -3667 348467
rect -3549 348349 240 348467
rect -4218 348338 240 348349
rect 291760 348627 296180 348638
rect 291760 348509 295511 348627
rect 295629 348509 296180 348627
rect 291760 348467 296180 348509
rect 291760 348349 295511 348467
rect 295629 348349 296180 348467
rect 291760 348338 296180 348349
rect -3758 348337 -3458 348338
rect 295420 348337 295720 348338
rect -2838 346838 -2538 346839
rect 294500 346838 294800 346839
rect -3298 346827 240 346838
rect -3298 346709 -2747 346827
rect -2629 346709 240 346827
rect -3298 346667 240 346709
rect -3298 346549 -2747 346667
rect -2629 346549 240 346667
rect -3298 346538 240 346549
rect 291760 346827 295260 346838
rect 291760 346709 294591 346827
rect 294709 346709 295260 346827
rect 291760 346667 295260 346709
rect 291760 346549 294591 346667
rect 294709 346549 295260 346667
rect 291760 346538 295260 346549
rect -2838 346537 -2538 346538
rect 294500 346537 294800 346538
rect -1918 345038 -1618 345039
rect 293580 345038 293880 345039
rect -2378 345027 240 345038
rect -2378 344909 -1827 345027
rect -1709 344909 240 345027
rect -2378 344867 240 344909
rect -2378 344749 -1827 344867
rect -1709 344749 240 344867
rect -2378 344738 240 344749
rect 291760 345027 294340 345038
rect 291760 344909 293671 345027
rect 293789 344909 294340 345027
rect 291760 344867 294340 344909
rect 291760 344749 293671 344867
rect 293789 344749 294340 344867
rect 291760 344738 294340 344749
rect -1918 344737 -1618 344738
rect 293580 344737 293880 344738
rect -998 343238 -698 343239
rect 292660 343238 292960 343239
rect -1458 343227 240 343238
rect -1458 343109 -907 343227
rect -789 343109 240 343227
rect -1458 343067 240 343109
rect -1458 342949 -907 343067
rect -789 342949 240 343067
rect -1458 342938 240 342949
rect 291760 343227 293420 343238
rect 291760 343109 292751 343227
rect 292869 343109 293420 343227
rect 291760 343067 293420 343109
rect 291760 342949 292751 343067
rect 292869 342949 293420 343067
rect 291760 342938 293420 342949
rect -998 342937 -698 342938
rect 292660 342937 292960 342938
rect -4218 339638 -3918 339639
rect 295880 339638 296180 339639
rect -4218 339627 240 339638
rect -4218 339509 -4127 339627
rect -4009 339509 240 339627
rect -4218 339467 240 339509
rect -4218 339349 -4127 339467
rect -4009 339349 240 339467
rect -4218 339338 240 339349
rect 291760 339627 296180 339638
rect 291760 339509 295971 339627
rect 296089 339509 296180 339627
rect 291760 339467 296180 339509
rect 291760 339349 295971 339467
rect 296089 339349 296180 339467
rect 291760 339338 296180 339349
rect -4218 339337 -3918 339338
rect 295880 339337 296180 339338
rect -3298 337838 -2998 337839
rect 294960 337838 295260 337839
rect -3298 337827 240 337838
rect -3298 337709 -3207 337827
rect -3089 337709 240 337827
rect -3298 337667 240 337709
rect -3298 337549 -3207 337667
rect -3089 337549 240 337667
rect -3298 337538 240 337549
rect 291760 337827 295260 337838
rect 291760 337709 295051 337827
rect 295169 337709 295260 337827
rect 291760 337667 295260 337709
rect 291760 337549 295051 337667
rect 295169 337549 295260 337667
rect 291760 337538 295260 337549
rect -3298 337537 -2998 337538
rect 294960 337537 295260 337538
rect -2378 336038 -2078 336039
rect 294040 336038 294340 336039
rect -2378 336027 240 336038
rect -2378 335909 -2287 336027
rect -2169 335909 240 336027
rect -2378 335867 240 335909
rect -2378 335749 -2287 335867
rect -2169 335749 240 335867
rect -2378 335738 240 335749
rect 291760 336027 294340 336038
rect 291760 335909 294131 336027
rect 294249 335909 294340 336027
rect 291760 335867 294340 335909
rect 291760 335749 294131 335867
rect 294249 335749 294340 335867
rect 291760 335738 294340 335749
rect -2378 335737 -2078 335738
rect 294040 335737 294340 335738
rect -1458 334238 -1158 334239
rect 293120 334238 293420 334239
rect -1458 334227 240 334238
rect -1458 334109 -1367 334227
rect -1249 334109 240 334227
rect -1458 334067 240 334109
rect -1458 333949 -1367 334067
rect -1249 333949 240 334067
rect -1458 333938 240 333949
rect 291760 334227 293420 334238
rect 291760 334109 293211 334227
rect 293329 334109 293420 334227
rect 291760 334067 293420 334109
rect 291760 333949 293211 334067
rect 293329 333949 293420 334067
rect 291760 333938 293420 333949
rect -1458 333937 -1158 333938
rect 293120 333937 293420 333938
rect -3758 330638 -3458 330639
rect 295420 330638 295720 330639
rect -4218 330627 240 330638
rect -4218 330509 -3667 330627
rect -3549 330509 240 330627
rect -4218 330467 240 330509
rect -4218 330349 -3667 330467
rect -3549 330349 240 330467
rect -4218 330338 240 330349
rect 291760 330627 296180 330638
rect 291760 330509 295511 330627
rect 295629 330509 296180 330627
rect 291760 330467 296180 330509
rect 291760 330349 295511 330467
rect 295629 330349 296180 330467
rect 291760 330338 296180 330349
rect -3758 330337 -3458 330338
rect 295420 330337 295720 330338
rect -2838 328838 -2538 328839
rect 294500 328838 294800 328839
rect -3298 328827 240 328838
rect -3298 328709 -2747 328827
rect -2629 328709 240 328827
rect -3298 328667 240 328709
rect -3298 328549 -2747 328667
rect -2629 328549 240 328667
rect -3298 328538 240 328549
rect 291760 328827 295260 328838
rect 291760 328709 294591 328827
rect 294709 328709 295260 328827
rect 291760 328667 295260 328709
rect 291760 328549 294591 328667
rect 294709 328549 295260 328667
rect 291760 328538 295260 328549
rect -2838 328537 -2538 328538
rect 294500 328537 294800 328538
rect -1918 327038 -1618 327039
rect 293580 327038 293880 327039
rect -2378 327027 240 327038
rect -2378 326909 -1827 327027
rect -1709 326909 240 327027
rect -2378 326867 240 326909
rect -2378 326749 -1827 326867
rect -1709 326749 240 326867
rect -2378 326738 240 326749
rect 291760 327027 294340 327038
rect 291760 326909 293671 327027
rect 293789 326909 294340 327027
rect 291760 326867 294340 326909
rect 291760 326749 293671 326867
rect 293789 326749 294340 326867
rect 291760 326738 294340 326749
rect -1918 326737 -1618 326738
rect 293580 326737 293880 326738
rect -998 325238 -698 325239
rect 292660 325238 292960 325239
rect -1458 325227 240 325238
rect -1458 325109 -907 325227
rect -789 325109 240 325227
rect -1458 325067 240 325109
rect -1458 324949 -907 325067
rect -789 324949 240 325067
rect -1458 324938 240 324949
rect 291760 325227 293420 325238
rect 291760 325109 292751 325227
rect 292869 325109 293420 325227
rect 291760 325067 293420 325109
rect 291760 324949 292751 325067
rect 292869 324949 293420 325067
rect 291760 324938 293420 324949
rect -998 324937 -698 324938
rect 292660 324937 292960 324938
rect -4218 321638 -3918 321639
rect 295880 321638 296180 321639
rect -4218 321627 240 321638
rect -4218 321509 -4127 321627
rect -4009 321509 240 321627
rect -4218 321467 240 321509
rect -4218 321349 -4127 321467
rect -4009 321349 240 321467
rect -4218 321338 240 321349
rect 291760 321627 296180 321638
rect 291760 321509 295971 321627
rect 296089 321509 296180 321627
rect 291760 321467 296180 321509
rect 291760 321349 295971 321467
rect 296089 321349 296180 321467
rect 291760 321338 296180 321349
rect -4218 321337 -3918 321338
rect 295880 321337 296180 321338
rect -3298 319838 -2998 319839
rect 294960 319838 295260 319839
rect -3298 319827 240 319838
rect -3298 319709 -3207 319827
rect -3089 319709 240 319827
rect -3298 319667 240 319709
rect -3298 319549 -3207 319667
rect -3089 319549 240 319667
rect -3298 319538 240 319549
rect 291760 319827 295260 319838
rect 291760 319709 295051 319827
rect 295169 319709 295260 319827
rect 291760 319667 295260 319709
rect 291760 319549 295051 319667
rect 295169 319549 295260 319667
rect 291760 319538 295260 319549
rect -3298 319537 -2998 319538
rect 294960 319537 295260 319538
rect -2378 318038 -2078 318039
rect 294040 318038 294340 318039
rect -2378 318027 240 318038
rect -2378 317909 -2287 318027
rect -2169 317909 240 318027
rect -2378 317867 240 317909
rect -2378 317749 -2287 317867
rect -2169 317749 240 317867
rect -2378 317738 240 317749
rect 291760 318027 294340 318038
rect 291760 317909 294131 318027
rect 294249 317909 294340 318027
rect 291760 317867 294340 317909
rect 291760 317749 294131 317867
rect 294249 317749 294340 317867
rect 291760 317738 294340 317749
rect -2378 317737 -2078 317738
rect 294040 317737 294340 317738
rect -1458 316238 -1158 316239
rect 293120 316238 293420 316239
rect -1458 316227 240 316238
rect -1458 316109 -1367 316227
rect -1249 316109 240 316227
rect -1458 316067 240 316109
rect -1458 315949 -1367 316067
rect -1249 315949 240 316067
rect -1458 315938 240 315949
rect 291760 316227 293420 316238
rect 291760 316109 293211 316227
rect 293329 316109 293420 316227
rect 291760 316067 293420 316109
rect 291760 315949 293211 316067
rect 293329 315949 293420 316067
rect 291760 315938 293420 315949
rect -1458 315937 -1158 315938
rect 293120 315937 293420 315938
rect -3758 312638 -3458 312639
rect 295420 312638 295720 312639
rect -4218 312627 240 312638
rect -4218 312509 -3667 312627
rect -3549 312509 240 312627
rect -4218 312467 240 312509
rect -4218 312349 -3667 312467
rect -3549 312349 240 312467
rect -4218 312338 240 312349
rect 291760 312627 296180 312638
rect 291760 312509 295511 312627
rect 295629 312509 296180 312627
rect 291760 312467 296180 312509
rect 291760 312349 295511 312467
rect 295629 312349 296180 312467
rect 291760 312338 296180 312349
rect -3758 312337 -3458 312338
rect 295420 312337 295720 312338
rect -2838 310838 -2538 310839
rect 294500 310838 294800 310839
rect -3298 310827 240 310838
rect -3298 310709 -2747 310827
rect -2629 310709 240 310827
rect -3298 310667 240 310709
rect -3298 310549 -2747 310667
rect -2629 310549 240 310667
rect -3298 310538 240 310549
rect 291760 310827 295260 310838
rect 291760 310709 294591 310827
rect 294709 310709 295260 310827
rect 291760 310667 295260 310709
rect 291760 310549 294591 310667
rect 294709 310549 295260 310667
rect 291760 310538 295260 310549
rect -2838 310537 -2538 310538
rect 294500 310537 294800 310538
rect -1918 309038 -1618 309039
rect 293580 309038 293880 309039
rect -2378 309027 240 309038
rect -2378 308909 -1827 309027
rect -1709 308909 240 309027
rect -2378 308867 240 308909
rect -2378 308749 -1827 308867
rect -1709 308749 240 308867
rect -2378 308738 240 308749
rect 291760 309027 294340 309038
rect 291760 308909 293671 309027
rect 293789 308909 294340 309027
rect 291760 308867 294340 308909
rect 291760 308749 293671 308867
rect 293789 308749 294340 308867
rect 291760 308738 294340 308749
rect -1918 308737 -1618 308738
rect 293580 308737 293880 308738
rect -998 307238 -698 307239
rect 292660 307238 292960 307239
rect -1458 307227 240 307238
rect -1458 307109 -907 307227
rect -789 307109 240 307227
rect -1458 307067 240 307109
rect -1458 306949 -907 307067
rect -789 306949 240 307067
rect -1458 306938 240 306949
rect 291760 307227 293420 307238
rect 291760 307109 292751 307227
rect 292869 307109 293420 307227
rect 291760 307067 293420 307109
rect 291760 306949 292751 307067
rect 292869 306949 293420 307067
rect 291760 306938 293420 306949
rect -998 306937 -698 306938
rect 292660 306937 292960 306938
rect -4218 303638 -3918 303639
rect 295880 303638 296180 303639
rect -4218 303627 240 303638
rect -4218 303509 -4127 303627
rect -4009 303509 240 303627
rect -4218 303467 240 303509
rect -4218 303349 -4127 303467
rect -4009 303349 240 303467
rect -4218 303338 240 303349
rect 291760 303627 296180 303638
rect 291760 303509 295971 303627
rect 296089 303509 296180 303627
rect 291760 303467 296180 303509
rect 291760 303349 295971 303467
rect 296089 303349 296180 303467
rect 291760 303338 296180 303349
rect -4218 303337 -3918 303338
rect 295880 303337 296180 303338
rect -3298 301838 -2998 301839
rect 294960 301838 295260 301839
rect -3298 301827 240 301838
rect -3298 301709 -3207 301827
rect -3089 301709 240 301827
rect -3298 301667 240 301709
rect -3298 301549 -3207 301667
rect -3089 301549 240 301667
rect -3298 301538 240 301549
rect 291760 301827 295260 301838
rect 291760 301709 295051 301827
rect 295169 301709 295260 301827
rect 291760 301667 295260 301709
rect 291760 301549 295051 301667
rect 295169 301549 295260 301667
rect 291760 301538 295260 301549
rect -3298 301537 -2998 301538
rect 294960 301537 295260 301538
rect -2378 300038 -2078 300039
rect 294040 300038 294340 300039
rect -2378 300027 240 300038
rect -2378 299909 -2287 300027
rect -2169 299909 240 300027
rect -2378 299867 240 299909
rect -2378 299749 -2287 299867
rect -2169 299749 240 299867
rect -2378 299738 240 299749
rect 291760 300027 294340 300038
rect 291760 299909 294131 300027
rect 294249 299909 294340 300027
rect 291760 299867 294340 299909
rect 291760 299749 294131 299867
rect 294249 299749 294340 299867
rect 291760 299738 294340 299749
rect -2378 299737 -2078 299738
rect 294040 299737 294340 299738
rect -1458 298238 -1158 298239
rect 293120 298238 293420 298239
rect -1458 298227 240 298238
rect -1458 298109 -1367 298227
rect -1249 298109 240 298227
rect -1458 298067 240 298109
rect -1458 297949 -1367 298067
rect -1249 297949 240 298067
rect -1458 297938 240 297949
rect 291760 298227 293420 298238
rect 291760 298109 293211 298227
rect 293329 298109 293420 298227
rect 291760 298067 293420 298109
rect 291760 297949 293211 298067
rect 293329 297949 293420 298067
rect 291760 297938 293420 297949
rect -1458 297937 -1158 297938
rect 293120 297937 293420 297938
rect -3758 294638 -3458 294639
rect 295420 294638 295720 294639
rect -4218 294627 240 294638
rect -4218 294509 -3667 294627
rect -3549 294509 240 294627
rect -4218 294467 240 294509
rect -4218 294349 -3667 294467
rect -3549 294349 240 294467
rect -4218 294338 240 294349
rect 291760 294627 296180 294638
rect 291760 294509 295511 294627
rect 295629 294509 296180 294627
rect 291760 294467 296180 294509
rect 291760 294349 295511 294467
rect 295629 294349 296180 294467
rect 291760 294338 296180 294349
rect -3758 294337 -3458 294338
rect 295420 294337 295720 294338
rect -2838 292838 -2538 292839
rect 294500 292838 294800 292839
rect -3298 292827 240 292838
rect -3298 292709 -2747 292827
rect -2629 292709 240 292827
rect -3298 292667 240 292709
rect -3298 292549 -2747 292667
rect -2629 292549 240 292667
rect -3298 292538 240 292549
rect 291760 292827 295260 292838
rect 291760 292709 294591 292827
rect 294709 292709 295260 292827
rect 291760 292667 295260 292709
rect 291760 292549 294591 292667
rect 294709 292549 295260 292667
rect 291760 292538 295260 292549
rect -2838 292537 -2538 292538
rect 294500 292537 294800 292538
rect -1918 291038 -1618 291039
rect 293580 291038 293880 291039
rect -2378 291027 240 291038
rect -2378 290909 -1827 291027
rect -1709 290909 240 291027
rect -2378 290867 240 290909
rect -2378 290749 -1827 290867
rect -1709 290749 240 290867
rect -2378 290738 240 290749
rect 291760 291027 294340 291038
rect 291760 290909 293671 291027
rect 293789 290909 294340 291027
rect 291760 290867 294340 290909
rect 291760 290749 293671 290867
rect 293789 290749 294340 290867
rect 291760 290738 294340 290749
rect -1918 290737 -1618 290738
rect 293580 290737 293880 290738
rect -998 289238 -698 289239
rect 292660 289238 292960 289239
rect -1458 289227 240 289238
rect -1458 289109 -907 289227
rect -789 289109 240 289227
rect -1458 289067 240 289109
rect -1458 288949 -907 289067
rect -789 288949 240 289067
rect -1458 288938 240 288949
rect 291760 289227 293420 289238
rect 291760 289109 292751 289227
rect 292869 289109 293420 289227
rect 291760 289067 293420 289109
rect 291760 288949 292751 289067
rect 292869 288949 293420 289067
rect 291760 288938 293420 288949
rect -998 288937 -698 288938
rect 292660 288937 292960 288938
rect -4218 285638 -3918 285639
rect 295880 285638 296180 285639
rect -4218 285627 240 285638
rect -4218 285509 -4127 285627
rect -4009 285509 240 285627
rect -4218 285467 240 285509
rect -4218 285349 -4127 285467
rect -4009 285349 240 285467
rect -4218 285338 240 285349
rect 291760 285627 296180 285638
rect 291760 285509 295971 285627
rect 296089 285509 296180 285627
rect 291760 285467 296180 285509
rect 291760 285349 295971 285467
rect 296089 285349 296180 285467
rect 291760 285338 296180 285349
rect -4218 285337 -3918 285338
rect 295880 285337 296180 285338
rect -3298 283838 -2998 283839
rect 294960 283838 295260 283839
rect -3298 283827 240 283838
rect -3298 283709 -3207 283827
rect -3089 283709 240 283827
rect -3298 283667 240 283709
rect -3298 283549 -3207 283667
rect -3089 283549 240 283667
rect -3298 283538 240 283549
rect 291760 283827 295260 283838
rect 291760 283709 295051 283827
rect 295169 283709 295260 283827
rect 291760 283667 295260 283709
rect 291760 283549 295051 283667
rect 295169 283549 295260 283667
rect 291760 283538 295260 283549
rect -3298 283537 -2998 283538
rect 294960 283537 295260 283538
rect -2378 282038 -2078 282039
rect 294040 282038 294340 282039
rect -2378 282027 240 282038
rect -2378 281909 -2287 282027
rect -2169 281909 240 282027
rect -2378 281867 240 281909
rect -2378 281749 -2287 281867
rect -2169 281749 240 281867
rect -2378 281738 240 281749
rect 291760 282027 294340 282038
rect 291760 281909 294131 282027
rect 294249 281909 294340 282027
rect 291760 281867 294340 281909
rect 291760 281749 294131 281867
rect 294249 281749 294340 281867
rect 291760 281738 294340 281749
rect -2378 281737 -2078 281738
rect 294040 281737 294340 281738
rect -1458 280238 -1158 280239
rect 293120 280238 293420 280239
rect -1458 280227 240 280238
rect -1458 280109 -1367 280227
rect -1249 280109 240 280227
rect -1458 280067 240 280109
rect -1458 279949 -1367 280067
rect -1249 279949 240 280067
rect -1458 279938 240 279949
rect 291760 280227 293420 280238
rect 291760 280109 293211 280227
rect 293329 280109 293420 280227
rect 291760 280067 293420 280109
rect 291760 279949 293211 280067
rect 293329 279949 293420 280067
rect 291760 279938 293420 279949
rect -1458 279937 -1158 279938
rect 293120 279937 293420 279938
rect -3758 276638 -3458 276639
rect 295420 276638 295720 276639
rect -4218 276627 240 276638
rect -4218 276509 -3667 276627
rect -3549 276509 240 276627
rect -4218 276467 240 276509
rect -4218 276349 -3667 276467
rect -3549 276349 240 276467
rect -4218 276338 240 276349
rect 291760 276627 296180 276638
rect 291760 276509 295511 276627
rect 295629 276509 296180 276627
rect 291760 276467 296180 276509
rect 291760 276349 295511 276467
rect 295629 276349 296180 276467
rect 291760 276338 296180 276349
rect -3758 276337 -3458 276338
rect 295420 276337 295720 276338
rect -2838 274838 -2538 274839
rect 294500 274838 294800 274839
rect -3298 274827 240 274838
rect -3298 274709 -2747 274827
rect -2629 274709 240 274827
rect -3298 274667 240 274709
rect -3298 274549 -2747 274667
rect -2629 274549 240 274667
rect -3298 274538 240 274549
rect 291760 274827 295260 274838
rect 291760 274709 294591 274827
rect 294709 274709 295260 274827
rect 291760 274667 295260 274709
rect 291760 274549 294591 274667
rect 294709 274549 295260 274667
rect 291760 274538 295260 274549
rect -2838 274537 -2538 274538
rect 294500 274537 294800 274538
rect -1918 273038 -1618 273039
rect 293580 273038 293880 273039
rect -2378 273027 240 273038
rect -2378 272909 -1827 273027
rect -1709 272909 240 273027
rect -2378 272867 240 272909
rect -2378 272749 -1827 272867
rect -1709 272749 240 272867
rect -2378 272738 240 272749
rect 291760 273027 294340 273038
rect 291760 272909 293671 273027
rect 293789 272909 294340 273027
rect 291760 272867 294340 272909
rect 291760 272749 293671 272867
rect 293789 272749 294340 272867
rect 291760 272738 294340 272749
rect -1918 272737 -1618 272738
rect 293580 272737 293880 272738
rect -998 271238 -698 271239
rect 292660 271238 292960 271239
rect -1458 271227 240 271238
rect -1458 271109 -907 271227
rect -789 271109 240 271227
rect -1458 271067 240 271109
rect -1458 270949 -907 271067
rect -789 270949 240 271067
rect -1458 270938 240 270949
rect 291760 271227 293420 271238
rect 291760 271109 292751 271227
rect 292869 271109 293420 271227
rect 291760 271067 293420 271109
rect 291760 270949 292751 271067
rect 292869 270949 293420 271067
rect 291760 270938 293420 270949
rect -998 270937 -698 270938
rect 292660 270937 292960 270938
rect -4218 267638 -3918 267639
rect 295880 267638 296180 267639
rect -4218 267627 240 267638
rect -4218 267509 -4127 267627
rect -4009 267509 240 267627
rect -4218 267467 240 267509
rect -4218 267349 -4127 267467
rect -4009 267349 240 267467
rect -4218 267338 240 267349
rect 291760 267627 296180 267638
rect 291760 267509 295971 267627
rect 296089 267509 296180 267627
rect 291760 267467 296180 267509
rect 291760 267349 295971 267467
rect 296089 267349 296180 267467
rect 291760 267338 296180 267349
rect -4218 267337 -3918 267338
rect 295880 267337 296180 267338
rect -3298 265838 -2998 265839
rect 294960 265838 295260 265839
rect -3298 265827 240 265838
rect -3298 265709 -3207 265827
rect -3089 265709 240 265827
rect -3298 265667 240 265709
rect -3298 265549 -3207 265667
rect -3089 265549 240 265667
rect -3298 265538 240 265549
rect 291760 265827 295260 265838
rect 291760 265709 295051 265827
rect 295169 265709 295260 265827
rect 291760 265667 295260 265709
rect 291760 265549 295051 265667
rect 295169 265549 295260 265667
rect 291760 265538 295260 265549
rect -3298 265537 -2998 265538
rect 294960 265537 295260 265538
rect -2378 264038 -2078 264039
rect 294040 264038 294340 264039
rect -2378 264027 240 264038
rect -2378 263909 -2287 264027
rect -2169 263909 240 264027
rect -2378 263867 240 263909
rect -2378 263749 -2287 263867
rect -2169 263749 240 263867
rect -2378 263738 240 263749
rect 291760 264027 294340 264038
rect 291760 263909 294131 264027
rect 294249 263909 294340 264027
rect 291760 263867 294340 263909
rect 291760 263749 294131 263867
rect 294249 263749 294340 263867
rect 291760 263738 294340 263749
rect -2378 263737 -2078 263738
rect 294040 263737 294340 263738
rect -1458 262238 -1158 262239
rect 293120 262238 293420 262239
rect -1458 262227 240 262238
rect -1458 262109 -1367 262227
rect -1249 262109 240 262227
rect -1458 262067 240 262109
rect -1458 261949 -1367 262067
rect -1249 261949 240 262067
rect -1458 261938 240 261949
rect 291760 262227 293420 262238
rect 291760 262109 293211 262227
rect 293329 262109 293420 262227
rect 291760 262067 293420 262109
rect 291760 261949 293211 262067
rect 293329 261949 293420 262067
rect 291760 261938 293420 261949
rect -1458 261937 -1158 261938
rect 293120 261937 293420 261938
rect -3758 258638 -3458 258639
rect 295420 258638 295720 258639
rect -4218 258627 240 258638
rect -4218 258509 -3667 258627
rect -3549 258509 240 258627
rect -4218 258467 240 258509
rect -4218 258349 -3667 258467
rect -3549 258349 240 258467
rect -4218 258338 240 258349
rect 291760 258627 296180 258638
rect 291760 258509 295511 258627
rect 295629 258509 296180 258627
rect 291760 258467 296180 258509
rect 291760 258349 295511 258467
rect 295629 258349 296180 258467
rect 291760 258338 296180 258349
rect -3758 258337 -3458 258338
rect 295420 258337 295720 258338
rect -2838 256838 -2538 256839
rect 294500 256838 294800 256839
rect -3298 256827 240 256838
rect -3298 256709 -2747 256827
rect -2629 256709 240 256827
rect -3298 256667 240 256709
rect -3298 256549 -2747 256667
rect -2629 256549 240 256667
rect -3298 256538 240 256549
rect 291760 256827 295260 256838
rect 291760 256709 294591 256827
rect 294709 256709 295260 256827
rect 291760 256667 295260 256709
rect 291760 256549 294591 256667
rect 294709 256549 295260 256667
rect 291760 256538 295260 256549
rect -2838 256537 -2538 256538
rect 294500 256537 294800 256538
rect -1918 255038 -1618 255039
rect 293580 255038 293880 255039
rect -2378 255027 240 255038
rect -2378 254909 -1827 255027
rect -1709 254909 240 255027
rect -2378 254867 240 254909
rect -2378 254749 -1827 254867
rect -1709 254749 240 254867
rect -2378 254738 240 254749
rect 291760 255027 294340 255038
rect 291760 254909 293671 255027
rect 293789 254909 294340 255027
rect 291760 254867 294340 254909
rect 291760 254749 293671 254867
rect 293789 254749 294340 254867
rect 291760 254738 294340 254749
rect -1918 254737 -1618 254738
rect 293580 254737 293880 254738
rect -998 253238 -698 253239
rect 292660 253238 292960 253239
rect -1458 253227 240 253238
rect -1458 253109 -907 253227
rect -789 253109 240 253227
rect -1458 253067 240 253109
rect -1458 252949 -907 253067
rect -789 252949 240 253067
rect -1458 252938 240 252949
rect 291760 253227 293420 253238
rect 291760 253109 292751 253227
rect 292869 253109 293420 253227
rect 291760 253067 293420 253109
rect 291760 252949 292751 253067
rect 292869 252949 293420 253067
rect 291760 252938 293420 252949
rect -998 252937 -698 252938
rect 292660 252937 292960 252938
rect -4218 249638 -3918 249639
rect 295880 249638 296180 249639
rect -4218 249627 240 249638
rect -4218 249509 -4127 249627
rect -4009 249509 240 249627
rect -4218 249467 240 249509
rect -4218 249349 -4127 249467
rect -4009 249349 240 249467
rect -4218 249338 240 249349
rect 291760 249627 296180 249638
rect 291760 249509 295971 249627
rect 296089 249509 296180 249627
rect 291760 249467 296180 249509
rect 291760 249349 295971 249467
rect 296089 249349 296180 249467
rect 291760 249338 296180 249349
rect -4218 249337 -3918 249338
rect 295880 249337 296180 249338
rect -3298 247838 -2998 247839
rect 294960 247838 295260 247839
rect -3298 247827 240 247838
rect -3298 247709 -3207 247827
rect -3089 247709 240 247827
rect -3298 247667 240 247709
rect -3298 247549 -3207 247667
rect -3089 247549 240 247667
rect -3298 247538 240 247549
rect 291760 247827 295260 247838
rect 291760 247709 295051 247827
rect 295169 247709 295260 247827
rect 291760 247667 295260 247709
rect 291760 247549 295051 247667
rect 295169 247549 295260 247667
rect 291760 247538 295260 247549
rect -3298 247537 -2998 247538
rect 294960 247537 295260 247538
rect -2378 246038 -2078 246039
rect 294040 246038 294340 246039
rect -2378 246027 240 246038
rect -2378 245909 -2287 246027
rect -2169 245909 240 246027
rect -2378 245867 240 245909
rect -2378 245749 -2287 245867
rect -2169 245749 240 245867
rect -2378 245738 240 245749
rect 291760 246027 294340 246038
rect 291760 245909 294131 246027
rect 294249 245909 294340 246027
rect 291760 245867 294340 245909
rect 291760 245749 294131 245867
rect 294249 245749 294340 245867
rect 291760 245738 294340 245749
rect -2378 245737 -2078 245738
rect 294040 245737 294340 245738
rect -1458 244238 -1158 244239
rect 293120 244238 293420 244239
rect -1458 244227 240 244238
rect -1458 244109 -1367 244227
rect -1249 244109 240 244227
rect -1458 244067 240 244109
rect -1458 243949 -1367 244067
rect -1249 243949 240 244067
rect -1458 243938 240 243949
rect 291760 244227 293420 244238
rect 291760 244109 293211 244227
rect 293329 244109 293420 244227
rect 291760 244067 293420 244109
rect 291760 243949 293211 244067
rect 293329 243949 293420 244067
rect 291760 243938 293420 243949
rect -1458 243937 -1158 243938
rect 293120 243937 293420 243938
rect -3758 240638 -3458 240639
rect 295420 240638 295720 240639
rect -4218 240627 240 240638
rect -4218 240509 -3667 240627
rect -3549 240509 240 240627
rect -4218 240467 240 240509
rect -4218 240349 -3667 240467
rect -3549 240349 240 240467
rect -4218 240338 240 240349
rect 291760 240627 296180 240638
rect 291760 240509 295511 240627
rect 295629 240509 296180 240627
rect 291760 240467 296180 240509
rect 291760 240349 295511 240467
rect 295629 240349 296180 240467
rect 291760 240338 296180 240349
rect -3758 240337 -3458 240338
rect 295420 240337 295720 240338
rect -2838 238838 -2538 238839
rect 294500 238838 294800 238839
rect -3298 238827 240 238838
rect -3298 238709 -2747 238827
rect -2629 238709 240 238827
rect -3298 238667 240 238709
rect -3298 238549 -2747 238667
rect -2629 238549 240 238667
rect -3298 238538 240 238549
rect 291760 238827 295260 238838
rect 291760 238709 294591 238827
rect 294709 238709 295260 238827
rect 291760 238667 295260 238709
rect 291760 238549 294591 238667
rect 294709 238549 295260 238667
rect 291760 238538 295260 238549
rect -2838 238537 -2538 238538
rect 294500 238537 294800 238538
rect -1918 237038 -1618 237039
rect 293580 237038 293880 237039
rect -2378 237027 240 237038
rect -2378 236909 -1827 237027
rect -1709 236909 240 237027
rect -2378 236867 240 236909
rect -2378 236749 -1827 236867
rect -1709 236749 240 236867
rect -2378 236738 240 236749
rect 291760 237027 294340 237038
rect 291760 236909 293671 237027
rect 293789 236909 294340 237027
rect 291760 236867 294340 236909
rect 291760 236749 293671 236867
rect 293789 236749 294340 236867
rect 291760 236738 294340 236749
rect -1918 236737 -1618 236738
rect 293580 236737 293880 236738
rect -998 235238 -698 235239
rect 292660 235238 292960 235239
rect -1458 235227 240 235238
rect -1458 235109 -907 235227
rect -789 235109 240 235227
rect -1458 235067 240 235109
rect -1458 234949 -907 235067
rect -789 234949 240 235067
rect -1458 234938 240 234949
rect 291760 235227 293420 235238
rect 291760 235109 292751 235227
rect 292869 235109 293420 235227
rect 291760 235067 293420 235109
rect 291760 234949 292751 235067
rect 292869 234949 293420 235067
rect 291760 234938 293420 234949
rect -998 234937 -698 234938
rect 292660 234937 292960 234938
rect -4218 231638 -3918 231639
rect 295880 231638 296180 231639
rect -4218 231627 240 231638
rect -4218 231509 -4127 231627
rect -4009 231509 240 231627
rect -4218 231467 240 231509
rect -4218 231349 -4127 231467
rect -4009 231349 240 231467
rect -4218 231338 240 231349
rect 291760 231627 296180 231638
rect 291760 231509 295971 231627
rect 296089 231509 296180 231627
rect 291760 231467 296180 231509
rect 291760 231349 295971 231467
rect 296089 231349 296180 231467
rect 291760 231338 296180 231349
rect -4218 231337 -3918 231338
rect 295880 231337 296180 231338
rect -3298 229838 -2998 229839
rect 294960 229838 295260 229839
rect -3298 229827 240 229838
rect -3298 229709 -3207 229827
rect -3089 229709 240 229827
rect -3298 229667 240 229709
rect -3298 229549 -3207 229667
rect -3089 229549 240 229667
rect -3298 229538 240 229549
rect 291760 229827 295260 229838
rect 291760 229709 295051 229827
rect 295169 229709 295260 229827
rect 291760 229667 295260 229709
rect 291760 229549 295051 229667
rect 295169 229549 295260 229667
rect 291760 229538 295260 229549
rect -3298 229537 -2998 229538
rect 294960 229537 295260 229538
rect -2378 228038 -2078 228039
rect 294040 228038 294340 228039
rect -2378 228027 240 228038
rect -2378 227909 -2287 228027
rect -2169 227909 240 228027
rect -2378 227867 240 227909
rect -2378 227749 -2287 227867
rect -2169 227749 240 227867
rect -2378 227738 240 227749
rect 291760 228027 294340 228038
rect 291760 227909 294131 228027
rect 294249 227909 294340 228027
rect 291760 227867 294340 227909
rect 291760 227749 294131 227867
rect 294249 227749 294340 227867
rect 291760 227738 294340 227749
rect -2378 227737 -2078 227738
rect 294040 227737 294340 227738
rect -1458 226238 -1158 226239
rect 293120 226238 293420 226239
rect -1458 226227 240 226238
rect -1458 226109 -1367 226227
rect -1249 226109 240 226227
rect -1458 226067 240 226109
rect -1458 225949 -1367 226067
rect -1249 225949 240 226067
rect -1458 225938 240 225949
rect 291760 226227 293420 226238
rect 291760 226109 293211 226227
rect 293329 226109 293420 226227
rect 291760 226067 293420 226109
rect 291760 225949 293211 226067
rect 293329 225949 293420 226067
rect 291760 225938 293420 225949
rect -1458 225937 -1158 225938
rect 293120 225937 293420 225938
rect -3758 222638 -3458 222639
rect 295420 222638 295720 222639
rect -4218 222627 240 222638
rect -4218 222509 -3667 222627
rect -3549 222509 240 222627
rect -4218 222467 240 222509
rect -4218 222349 -3667 222467
rect -3549 222349 240 222467
rect -4218 222338 240 222349
rect 291760 222627 296180 222638
rect 291760 222509 295511 222627
rect 295629 222509 296180 222627
rect 291760 222467 296180 222509
rect 291760 222349 295511 222467
rect 295629 222349 296180 222467
rect 291760 222338 296180 222349
rect -3758 222337 -3458 222338
rect 295420 222337 295720 222338
rect -2838 220838 -2538 220839
rect 294500 220838 294800 220839
rect -3298 220827 240 220838
rect -3298 220709 -2747 220827
rect -2629 220709 240 220827
rect -3298 220667 240 220709
rect -3298 220549 -2747 220667
rect -2629 220549 240 220667
rect -3298 220538 240 220549
rect 291760 220827 295260 220838
rect 291760 220709 294591 220827
rect 294709 220709 295260 220827
rect 291760 220667 295260 220709
rect 291760 220549 294591 220667
rect 294709 220549 295260 220667
rect 291760 220538 295260 220549
rect -2838 220537 -2538 220538
rect 294500 220537 294800 220538
rect -1918 219038 -1618 219039
rect 293580 219038 293880 219039
rect -2378 219027 240 219038
rect -2378 218909 -1827 219027
rect -1709 218909 240 219027
rect -2378 218867 240 218909
rect -2378 218749 -1827 218867
rect -1709 218749 240 218867
rect -2378 218738 240 218749
rect 291760 219027 294340 219038
rect 291760 218909 293671 219027
rect 293789 218909 294340 219027
rect 291760 218867 294340 218909
rect 291760 218749 293671 218867
rect 293789 218749 294340 218867
rect 291760 218738 294340 218749
rect -1918 218737 -1618 218738
rect 293580 218737 293880 218738
rect -998 217238 -698 217239
rect 292660 217238 292960 217239
rect -1458 217227 240 217238
rect -1458 217109 -907 217227
rect -789 217109 240 217227
rect -1458 217067 240 217109
rect -1458 216949 -907 217067
rect -789 216949 240 217067
rect -1458 216938 240 216949
rect 291760 217227 293420 217238
rect 291760 217109 292751 217227
rect 292869 217109 293420 217227
rect 291760 217067 293420 217109
rect 291760 216949 292751 217067
rect 292869 216949 293420 217067
rect 291760 216938 293420 216949
rect -998 216937 -698 216938
rect 292660 216937 292960 216938
rect -4218 213638 -3918 213639
rect 295880 213638 296180 213639
rect -4218 213627 240 213638
rect -4218 213509 -4127 213627
rect -4009 213509 240 213627
rect -4218 213467 240 213509
rect -4218 213349 -4127 213467
rect -4009 213349 240 213467
rect -4218 213338 240 213349
rect 291760 213627 296180 213638
rect 291760 213509 295971 213627
rect 296089 213509 296180 213627
rect 291760 213467 296180 213509
rect 291760 213349 295971 213467
rect 296089 213349 296180 213467
rect 291760 213338 296180 213349
rect -4218 213337 -3918 213338
rect 295880 213337 296180 213338
rect -3298 211838 -2998 211839
rect 294960 211838 295260 211839
rect -3298 211827 240 211838
rect -3298 211709 -3207 211827
rect -3089 211709 240 211827
rect -3298 211667 240 211709
rect -3298 211549 -3207 211667
rect -3089 211549 240 211667
rect -3298 211538 240 211549
rect 291760 211827 295260 211838
rect 291760 211709 295051 211827
rect 295169 211709 295260 211827
rect 291760 211667 295260 211709
rect 291760 211549 295051 211667
rect 295169 211549 295260 211667
rect 291760 211538 295260 211549
rect -3298 211537 -2998 211538
rect 294960 211537 295260 211538
rect -2378 210038 -2078 210039
rect 294040 210038 294340 210039
rect -2378 210027 240 210038
rect -2378 209909 -2287 210027
rect -2169 209909 240 210027
rect -2378 209867 240 209909
rect -2378 209749 -2287 209867
rect -2169 209749 240 209867
rect -2378 209738 240 209749
rect 291760 210027 294340 210038
rect 291760 209909 294131 210027
rect 294249 209909 294340 210027
rect 291760 209867 294340 209909
rect 291760 209749 294131 209867
rect 294249 209749 294340 209867
rect 291760 209738 294340 209749
rect -2378 209737 -2078 209738
rect 294040 209737 294340 209738
rect -1458 208238 -1158 208239
rect 293120 208238 293420 208239
rect -1458 208227 240 208238
rect -1458 208109 -1367 208227
rect -1249 208109 240 208227
rect -1458 208067 240 208109
rect -1458 207949 -1367 208067
rect -1249 207949 240 208067
rect -1458 207938 240 207949
rect 291760 208227 293420 208238
rect 291760 208109 293211 208227
rect 293329 208109 293420 208227
rect 291760 208067 293420 208109
rect 291760 207949 293211 208067
rect 293329 207949 293420 208067
rect 291760 207938 293420 207949
rect -1458 207937 -1158 207938
rect 293120 207937 293420 207938
rect -3758 204638 -3458 204639
rect 295420 204638 295720 204639
rect -4218 204627 240 204638
rect -4218 204509 -3667 204627
rect -3549 204509 240 204627
rect -4218 204467 240 204509
rect -4218 204349 -3667 204467
rect -3549 204349 240 204467
rect -4218 204338 240 204349
rect 291760 204627 296180 204638
rect 291760 204509 295511 204627
rect 295629 204509 296180 204627
rect 291760 204467 296180 204509
rect 291760 204349 295511 204467
rect 295629 204349 296180 204467
rect 291760 204338 296180 204349
rect -3758 204337 -3458 204338
rect 295420 204337 295720 204338
rect -2838 202838 -2538 202839
rect 294500 202838 294800 202839
rect -3298 202827 240 202838
rect -3298 202709 -2747 202827
rect -2629 202709 240 202827
rect -3298 202667 240 202709
rect -3298 202549 -2747 202667
rect -2629 202549 240 202667
rect -3298 202538 240 202549
rect 291760 202827 295260 202838
rect 291760 202709 294591 202827
rect 294709 202709 295260 202827
rect 291760 202667 295260 202709
rect 291760 202549 294591 202667
rect 294709 202549 295260 202667
rect 291760 202538 295260 202549
rect -2838 202537 -2538 202538
rect 294500 202537 294800 202538
rect -1918 201038 -1618 201039
rect 293580 201038 293880 201039
rect -2378 201027 240 201038
rect -2378 200909 -1827 201027
rect -1709 200909 240 201027
rect -2378 200867 240 200909
rect -2378 200749 -1827 200867
rect -1709 200749 240 200867
rect -2378 200738 240 200749
rect 291760 201027 294340 201038
rect 291760 200909 293671 201027
rect 293789 200909 294340 201027
rect 291760 200867 294340 200909
rect 291760 200749 293671 200867
rect 293789 200749 294340 200867
rect 291760 200738 294340 200749
rect -1918 200737 -1618 200738
rect 293580 200737 293880 200738
rect -998 199238 -698 199239
rect 292660 199238 292960 199239
rect -1458 199227 240 199238
rect -1458 199109 -907 199227
rect -789 199109 240 199227
rect -1458 199067 240 199109
rect -1458 198949 -907 199067
rect -789 198949 240 199067
rect -1458 198938 240 198949
rect 291760 199227 293420 199238
rect 291760 199109 292751 199227
rect 292869 199109 293420 199227
rect 291760 199067 293420 199109
rect 291760 198949 292751 199067
rect 292869 198949 293420 199067
rect 291760 198938 293420 198949
rect -998 198937 -698 198938
rect 292660 198937 292960 198938
rect -4218 195638 -3918 195639
rect 295880 195638 296180 195639
rect -4218 195627 240 195638
rect -4218 195509 -4127 195627
rect -4009 195509 240 195627
rect -4218 195467 240 195509
rect -4218 195349 -4127 195467
rect -4009 195349 240 195467
rect -4218 195338 240 195349
rect 291760 195627 296180 195638
rect 291760 195509 295971 195627
rect 296089 195509 296180 195627
rect 291760 195467 296180 195509
rect 291760 195349 295971 195467
rect 296089 195349 296180 195467
rect 291760 195338 296180 195349
rect -4218 195337 -3918 195338
rect 295880 195337 296180 195338
rect -3298 193838 -2998 193839
rect 294960 193838 295260 193839
rect -3298 193827 240 193838
rect -3298 193709 -3207 193827
rect -3089 193709 240 193827
rect -3298 193667 240 193709
rect -3298 193549 -3207 193667
rect -3089 193549 240 193667
rect -3298 193538 240 193549
rect 291760 193827 295260 193838
rect 291760 193709 295051 193827
rect 295169 193709 295260 193827
rect 291760 193667 295260 193709
rect 291760 193549 295051 193667
rect 295169 193549 295260 193667
rect 291760 193538 295260 193549
rect -3298 193537 -2998 193538
rect 294960 193537 295260 193538
rect -2378 192038 -2078 192039
rect 294040 192038 294340 192039
rect -2378 192027 240 192038
rect -2378 191909 -2287 192027
rect -2169 191909 240 192027
rect -2378 191867 240 191909
rect -2378 191749 -2287 191867
rect -2169 191749 240 191867
rect -2378 191738 240 191749
rect 291760 192027 294340 192038
rect 291760 191909 294131 192027
rect 294249 191909 294340 192027
rect 291760 191867 294340 191909
rect 291760 191749 294131 191867
rect 294249 191749 294340 191867
rect 291760 191738 294340 191749
rect -2378 191737 -2078 191738
rect 294040 191737 294340 191738
rect -1458 190238 -1158 190239
rect 293120 190238 293420 190239
rect -1458 190227 240 190238
rect -1458 190109 -1367 190227
rect -1249 190109 240 190227
rect -1458 190067 240 190109
rect -1458 189949 -1367 190067
rect -1249 189949 240 190067
rect -1458 189938 240 189949
rect 291760 190227 293420 190238
rect 291760 190109 293211 190227
rect 293329 190109 293420 190227
rect 291760 190067 293420 190109
rect 291760 189949 293211 190067
rect 293329 189949 293420 190067
rect 291760 189938 293420 189949
rect -1458 189937 -1158 189938
rect 293120 189937 293420 189938
rect -3758 186638 -3458 186639
rect 295420 186638 295720 186639
rect -4218 186627 240 186638
rect -4218 186509 -3667 186627
rect -3549 186509 240 186627
rect -4218 186467 240 186509
rect -4218 186349 -3667 186467
rect -3549 186349 240 186467
rect -4218 186338 240 186349
rect 291760 186627 296180 186638
rect 291760 186509 295511 186627
rect 295629 186509 296180 186627
rect 291760 186467 296180 186509
rect 291760 186349 295511 186467
rect 295629 186349 296180 186467
rect 291760 186338 296180 186349
rect -3758 186337 -3458 186338
rect 295420 186337 295720 186338
rect -2838 184838 -2538 184839
rect 294500 184838 294800 184839
rect -3298 184827 240 184838
rect -3298 184709 -2747 184827
rect -2629 184709 240 184827
rect -3298 184667 240 184709
rect -3298 184549 -2747 184667
rect -2629 184549 240 184667
rect -3298 184538 240 184549
rect 291760 184827 295260 184838
rect 291760 184709 294591 184827
rect 294709 184709 295260 184827
rect 291760 184667 295260 184709
rect 291760 184549 294591 184667
rect 294709 184549 295260 184667
rect 291760 184538 295260 184549
rect -2838 184537 -2538 184538
rect 294500 184537 294800 184538
rect -1918 183038 -1618 183039
rect 293580 183038 293880 183039
rect -2378 183027 240 183038
rect -2378 182909 -1827 183027
rect -1709 182909 240 183027
rect -2378 182867 240 182909
rect -2378 182749 -1827 182867
rect -1709 182749 240 182867
rect -2378 182738 240 182749
rect 291760 183027 294340 183038
rect 291760 182909 293671 183027
rect 293789 182909 294340 183027
rect 291760 182867 294340 182909
rect 291760 182749 293671 182867
rect 293789 182749 294340 182867
rect 291760 182738 294340 182749
rect -1918 182737 -1618 182738
rect 293580 182737 293880 182738
rect -998 181238 -698 181239
rect 292660 181238 292960 181239
rect -1458 181227 240 181238
rect -1458 181109 -907 181227
rect -789 181109 240 181227
rect -1458 181067 240 181109
rect -1458 180949 -907 181067
rect -789 180949 240 181067
rect -1458 180938 240 180949
rect 291760 181227 293420 181238
rect 291760 181109 292751 181227
rect 292869 181109 293420 181227
rect 291760 181067 293420 181109
rect 291760 180949 292751 181067
rect 292869 180949 293420 181067
rect 291760 180938 293420 180949
rect -998 180937 -698 180938
rect 292660 180937 292960 180938
rect -4218 177638 -3918 177639
rect 295880 177638 296180 177639
rect -4218 177627 240 177638
rect -4218 177509 -4127 177627
rect -4009 177509 240 177627
rect -4218 177467 240 177509
rect -4218 177349 -4127 177467
rect -4009 177349 240 177467
rect -4218 177338 240 177349
rect 291760 177627 296180 177638
rect 291760 177509 295971 177627
rect 296089 177509 296180 177627
rect 291760 177467 296180 177509
rect 291760 177349 295971 177467
rect 296089 177349 296180 177467
rect 291760 177338 296180 177349
rect -4218 177337 -3918 177338
rect 295880 177337 296180 177338
rect -3298 175838 -2998 175839
rect 294960 175838 295260 175839
rect -3298 175827 240 175838
rect -3298 175709 -3207 175827
rect -3089 175709 240 175827
rect -3298 175667 240 175709
rect -3298 175549 -3207 175667
rect -3089 175549 240 175667
rect -3298 175538 240 175549
rect 291760 175827 295260 175838
rect 291760 175709 295051 175827
rect 295169 175709 295260 175827
rect 291760 175667 295260 175709
rect 291760 175549 295051 175667
rect 295169 175549 295260 175667
rect 291760 175538 295260 175549
rect -3298 175537 -2998 175538
rect 294960 175537 295260 175538
rect -2378 174038 -2078 174039
rect 294040 174038 294340 174039
rect -2378 174027 240 174038
rect -2378 173909 -2287 174027
rect -2169 173909 240 174027
rect -2378 173867 240 173909
rect -2378 173749 -2287 173867
rect -2169 173749 240 173867
rect -2378 173738 240 173749
rect 291760 174027 294340 174038
rect 291760 173909 294131 174027
rect 294249 173909 294340 174027
rect 291760 173867 294340 173909
rect 291760 173749 294131 173867
rect 294249 173749 294340 173867
rect 291760 173738 294340 173749
rect -2378 173737 -2078 173738
rect 294040 173737 294340 173738
rect -1458 172238 -1158 172239
rect 293120 172238 293420 172239
rect -1458 172227 240 172238
rect -1458 172109 -1367 172227
rect -1249 172109 240 172227
rect -1458 172067 240 172109
rect -1458 171949 -1367 172067
rect -1249 171949 240 172067
rect -1458 171938 240 171949
rect 291760 172227 293420 172238
rect 291760 172109 293211 172227
rect 293329 172109 293420 172227
rect 291760 172067 293420 172109
rect 291760 171949 293211 172067
rect 293329 171949 293420 172067
rect 291760 171938 293420 171949
rect -1458 171937 -1158 171938
rect 293120 171937 293420 171938
rect -3758 168638 -3458 168639
rect 295420 168638 295720 168639
rect -4218 168627 240 168638
rect -4218 168509 -3667 168627
rect -3549 168509 240 168627
rect -4218 168467 240 168509
rect -4218 168349 -3667 168467
rect -3549 168349 240 168467
rect -4218 168338 240 168349
rect 291760 168627 296180 168638
rect 291760 168509 295511 168627
rect 295629 168509 296180 168627
rect 291760 168467 296180 168509
rect 291760 168349 295511 168467
rect 295629 168349 296180 168467
rect 291760 168338 296180 168349
rect -3758 168337 -3458 168338
rect 295420 168337 295720 168338
rect -2838 166838 -2538 166839
rect 294500 166838 294800 166839
rect -3298 166827 240 166838
rect -3298 166709 -2747 166827
rect -2629 166709 240 166827
rect -3298 166667 240 166709
rect -3298 166549 -2747 166667
rect -2629 166549 240 166667
rect -3298 166538 240 166549
rect 291760 166827 295260 166838
rect 291760 166709 294591 166827
rect 294709 166709 295260 166827
rect 291760 166667 295260 166709
rect 291760 166549 294591 166667
rect 294709 166549 295260 166667
rect 291760 166538 295260 166549
rect -2838 166537 -2538 166538
rect 294500 166537 294800 166538
rect -1918 165038 -1618 165039
rect 293580 165038 293880 165039
rect -2378 165027 240 165038
rect -2378 164909 -1827 165027
rect -1709 164909 240 165027
rect -2378 164867 240 164909
rect -2378 164749 -1827 164867
rect -1709 164749 240 164867
rect -2378 164738 240 164749
rect 291760 165027 294340 165038
rect 291760 164909 293671 165027
rect 293789 164909 294340 165027
rect 291760 164867 294340 164909
rect 291760 164749 293671 164867
rect 293789 164749 294340 164867
rect 291760 164738 294340 164749
rect -1918 164737 -1618 164738
rect 293580 164737 293880 164738
rect -998 163238 -698 163239
rect 292660 163238 292960 163239
rect -1458 163227 240 163238
rect -1458 163109 -907 163227
rect -789 163109 240 163227
rect -1458 163067 240 163109
rect -1458 162949 -907 163067
rect -789 162949 240 163067
rect -1458 162938 240 162949
rect 291760 163227 293420 163238
rect 291760 163109 292751 163227
rect 292869 163109 293420 163227
rect 291760 163067 293420 163109
rect 291760 162949 292751 163067
rect 292869 162949 293420 163067
rect 291760 162938 293420 162949
rect -998 162937 -698 162938
rect 292660 162937 292960 162938
rect -4218 159638 -3918 159639
rect 295880 159638 296180 159639
rect -4218 159627 240 159638
rect -4218 159509 -4127 159627
rect -4009 159509 240 159627
rect -4218 159467 240 159509
rect -4218 159349 -4127 159467
rect -4009 159349 240 159467
rect -4218 159338 240 159349
rect 291760 159627 296180 159638
rect 291760 159509 295971 159627
rect 296089 159509 296180 159627
rect 291760 159467 296180 159509
rect 291760 159349 295971 159467
rect 296089 159349 296180 159467
rect 291760 159338 296180 159349
rect -4218 159337 -3918 159338
rect 295880 159337 296180 159338
rect -3298 157838 -2998 157839
rect 294960 157838 295260 157839
rect -3298 157827 240 157838
rect -3298 157709 -3207 157827
rect -3089 157709 240 157827
rect -3298 157667 240 157709
rect -3298 157549 -3207 157667
rect -3089 157549 240 157667
rect -3298 157538 240 157549
rect 291760 157827 295260 157838
rect 291760 157709 295051 157827
rect 295169 157709 295260 157827
rect 291760 157667 295260 157709
rect 291760 157549 295051 157667
rect 295169 157549 295260 157667
rect 291760 157538 295260 157549
rect -3298 157537 -2998 157538
rect 294960 157537 295260 157538
rect -2378 156038 -2078 156039
rect 294040 156038 294340 156039
rect -2378 156027 240 156038
rect -2378 155909 -2287 156027
rect -2169 155909 240 156027
rect -2378 155867 240 155909
rect -2378 155749 -2287 155867
rect -2169 155749 240 155867
rect -2378 155738 240 155749
rect 291760 156027 294340 156038
rect 291760 155909 294131 156027
rect 294249 155909 294340 156027
rect 291760 155867 294340 155909
rect 291760 155749 294131 155867
rect 294249 155749 294340 155867
rect 291760 155738 294340 155749
rect -2378 155737 -2078 155738
rect 294040 155737 294340 155738
rect -1458 154238 -1158 154239
rect 293120 154238 293420 154239
rect -1458 154227 240 154238
rect -1458 154109 -1367 154227
rect -1249 154109 240 154227
rect -1458 154067 240 154109
rect -1458 153949 -1367 154067
rect -1249 153949 240 154067
rect -1458 153938 240 153949
rect 291760 154227 293420 154238
rect 291760 154109 293211 154227
rect 293329 154109 293420 154227
rect 291760 154067 293420 154109
rect 291760 153949 293211 154067
rect 293329 153949 293420 154067
rect 291760 153938 293420 153949
rect -1458 153937 -1158 153938
rect 293120 153937 293420 153938
rect -3758 150638 -3458 150639
rect 295420 150638 295720 150639
rect -4218 150627 240 150638
rect -4218 150509 -3667 150627
rect -3549 150509 240 150627
rect -4218 150467 240 150509
rect -4218 150349 -3667 150467
rect -3549 150349 240 150467
rect -4218 150338 240 150349
rect 291760 150627 296180 150638
rect 291760 150509 295511 150627
rect 295629 150509 296180 150627
rect 291760 150467 296180 150509
rect 291760 150349 295511 150467
rect 295629 150349 296180 150467
rect 291760 150338 296180 150349
rect -3758 150337 -3458 150338
rect 295420 150337 295720 150338
rect -2838 148838 -2538 148839
rect 294500 148838 294800 148839
rect -3298 148827 240 148838
rect -3298 148709 -2747 148827
rect -2629 148709 240 148827
rect -3298 148667 240 148709
rect -3298 148549 -2747 148667
rect -2629 148549 240 148667
rect -3298 148538 240 148549
rect 291760 148827 295260 148838
rect 291760 148709 294591 148827
rect 294709 148709 295260 148827
rect 291760 148667 295260 148709
rect 291760 148549 294591 148667
rect 294709 148549 295260 148667
rect 291760 148538 295260 148549
rect -2838 148537 -2538 148538
rect 294500 148537 294800 148538
rect -1918 147038 -1618 147039
rect 293580 147038 293880 147039
rect -2378 147027 240 147038
rect -2378 146909 -1827 147027
rect -1709 146909 240 147027
rect -2378 146867 240 146909
rect -2378 146749 -1827 146867
rect -1709 146749 240 146867
rect -2378 146738 240 146749
rect 291760 147027 294340 147038
rect 291760 146909 293671 147027
rect 293789 146909 294340 147027
rect 291760 146867 294340 146909
rect 291760 146749 293671 146867
rect 293789 146749 294340 146867
rect 291760 146738 294340 146749
rect -1918 146737 -1618 146738
rect 293580 146737 293880 146738
rect -998 145238 -698 145239
rect 292660 145238 292960 145239
rect -1458 145227 240 145238
rect -1458 145109 -907 145227
rect -789 145109 240 145227
rect -1458 145067 240 145109
rect -1458 144949 -907 145067
rect -789 144949 240 145067
rect -1458 144938 240 144949
rect 291760 145227 293420 145238
rect 291760 145109 292751 145227
rect 292869 145109 293420 145227
rect 291760 145067 293420 145109
rect 291760 144949 292751 145067
rect 292869 144949 293420 145067
rect 291760 144938 293420 144949
rect -998 144937 -698 144938
rect 292660 144937 292960 144938
rect -4218 141638 -3918 141639
rect 295880 141638 296180 141639
rect -4218 141627 240 141638
rect -4218 141509 -4127 141627
rect -4009 141509 240 141627
rect -4218 141467 240 141509
rect -4218 141349 -4127 141467
rect -4009 141349 240 141467
rect -4218 141338 240 141349
rect 291760 141627 296180 141638
rect 291760 141509 295971 141627
rect 296089 141509 296180 141627
rect 291760 141467 296180 141509
rect 291760 141349 295971 141467
rect 296089 141349 296180 141467
rect 291760 141338 296180 141349
rect -4218 141337 -3918 141338
rect 295880 141337 296180 141338
rect -3298 139838 -2998 139839
rect 294960 139838 295260 139839
rect -3298 139827 240 139838
rect -3298 139709 -3207 139827
rect -3089 139709 240 139827
rect -3298 139667 240 139709
rect -3298 139549 -3207 139667
rect -3089 139549 240 139667
rect -3298 139538 240 139549
rect 291760 139827 295260 139838
rect 291760 139709 295051 139827
rect 295169 139709 295260 139827
rect 291760 139667 295260 139709
rect 291760 139549 295051 139667
rect 295169 139549 295260 139667
rect 291760 139538 295260 139549
rect -3298 139537 -2998 139538
rect 294960 139537 295260 139538
rect -2378 138038 -2078 138039
rect 294040 138038 294340 138039
rect -2378 138027 240 138038
rect -2378 137909 -2287 138027
rect -2169 137909 240 138027
rect -2378 137867 240 137909
rect -2378 137749 -2287 137867
rect -2169 137749 240 137867
rect -2378 137738 240 137749
rect 291760 138027 294340 138038
rect 291760 137909 294131 138027
rect 294249 137909 294340 138027
rect 291760 137867 294340 137909
rect 291760 137749 294131 137867
rect 294249 137749 294340 137867
rect 291760 137738 294340 137749
rect -2378 137737 -2078 137738
rect 294040 137737 294340 137738
rect -1458 136238 -1158 136239
rect 293120 136238 293420 136239
rect -1458 136227 240 136238
rect -1458 136109 -1367 136227
rect -1249 136109 240 136227
rect -1458 136067 240 136109
rect -1458 135949 -1367 136067
rect -1249 135949 240 136067
rect -1458 135938 240 135949
rect 291760 136227 293420 136238
rect 291760 136109 293211 136227
rect 293329 136109 293420 136227
rect 291760 136067 293420 136109
rect 291760 135949 293211 136067
rect 293329 135949 293420 136067
rect 291760 135938 293420 135949
rect -1458 135937 -1158 135938
rect 293120 135937 293420 135938
rect -3758 132638 -3458 132639
rect 295420 132638 295720 132639
rect -4218 132627 240 132638
rect -4218 132509 -3667 132627
rect -3549 132509 240 132627
rect -4218 132467 240 132509
rect -4218 132349 -3667 132467
rect -3549 132349 240 132467
rect -4218 132338 240 132349
rect 291760 132627 296180 132638
rect 291760 132509 295511 132627
rect 295629 132509 296180 132627
rect 291760 132467 296180 132509
rect 291760 132349 295511 132467
rect 295629 132349 296180 132467
rect 291760 132338 296180 132349
rect -3758 132337 -3458 132338
rect 295420 132337 295720 132338
rect -2838 130838 -2538 130839
rect 294500 130838 294800 130839
rect -3298 130827 240 130838
rect -3298 130709 -2747 130827
rect -2629 130709 240 130827
rect -3298 130667 240 130709
rect -3298 130549 -2747 130667
rect -2629 130549 240 130667
rect -3298 130538 240 130549
rect 291760 130827 295260 130838
rect 291760 130709 294591 130827
rect 294709 130709 295260 130827
rect 291760 130667 295260 130709
rect 291760 130549 294591 130667
rect 294709 130549 295260 130667
rect 291760 130538 295260 130549
rect -2838 130537 -2538 130538
rect 294500 130537 294800 130538
rect -1918 129038 -1618 129039
rect 293580 129038 293880 129039
rect -2378 129027 240 129038
rect -2378 128909 -1827 129027
rect -1709 128909 240 129027
rect -2378 128867 240 128909
rect -2378 128749 -1827 128867
rect -1709 128749 240 128867
rect -2378 128738 240 128749
rect 291760 129027 294340 129038
rect 291760 128909 293671 129027
rect 293789 128909 294340 129027
rect 291760 128867 294340 128909
rect 291760 128749 293671 128867
rect 293789 128749 294340 128867
rect 291760 128738 294340 128749
rect -1918 128737 -1618 128738
rect 293580 128737 293880 128738
rect -998 127238 -698 127239
rect 292660 127238 292960 127239
rect -1458 127227 240 127238
rect -1458 127109 -907 127227
rect -789 127109 240 127227
rect -1458 127067 240 127109
rect -1458 126949 -907 127067
rect -789 126949 240 127067
rect -1458 126938 240 126949
rect 291760 127227 293420 127238
rect 291760 127109 292751 127227
rect 292869 127109 293420 127227
rect 291760 127067 293420 127109
rect 291760 126949 292751 127067
rect 292869 126949 293420 127067
rect 291760 126938 293420 126949
rect -998 126937 -698 126938
rect 292660 126937 292960 126938
rect -4218 123638 -3918 123639
rect 295880 123638 296180 123639
rect -4218 123627 240 123638
rect -4218 123509 -4127 123627
rect -4009 123509 240 123627
rect -4218 123467 240 123509
rect -4218 123349 -4127 123467
rect -4009 123349 240 123467
rect -4218 123338 240 123349
rect 291760 123627 296180 123638
rect 291760 123509 295971 123627
rect 296089 123509 296180 123627
rect 291760 123467 296180 123509
rect 291760 123349 295971 123467
rect 296089 123349 296180 123467
rect 291760 123338 296180 123349
rect -4218 123337 -3918 123338
rect 295880 123337 296180 123338
rect -3298 121838 -2998 121839
rect 294960 121838 295260 121839
rect -3298 121827 240 121838
rect -3298 121709 -3207 121827
rect -3089 121709 240 121827
rect -3298 121667 240 121709
rect -3298 121549 -3207 121667
rect -3089 121549 240 121667
rect -3298 121538 240 121549
rect 291760 121827 295260 121838
rect 291760 121709 295051 121827
rect 295169 121709 295260 121827
rect 291760 121667 295260 121709
rect 291760 121549 295051 121667
rect 295169 121549 295260 121667
rect 291760 121538 295260 121549
rect -3298 121537 -2998 121538
rect 294960 121537 295260 121538
rect -2378 120038 -2078 120039
rect 294040 120038 294340 120039
rect -2378 120027 240 120038
rect -2378 119909 -2287 120027
rect -2169 119909 240 120027
rect -2378 119867 240 119909
rect -2378 119749 -2287 119867
rect -2169 119749 240 119867
rect -2378 119738 240 119749
rect 291760 120027 294340 120038
rect 291760 119909 294131 120027
rect 294249 119909 294340 120027
rect 291760 119867 294340 119909
rect 291760 119749 294131 119867
rect 294249 119749 294340 119867
rect 291760 119738 294340 119749
rect -2378 119737 -2078 119738
rect 294040 119737 294340 119738
rect -1458 118238 -1158 118239
rect 293120 118238 293420 118239
rect -1458 118227 240 118238
rect -1458 118109 -1367 118227
rect -1249 118109 240 118227
rect -1458 118067 240 118109
rect -1458 117949 -1367 118067
rect -1249 117949 240 118067
rect -1458 117938 240 117949
rect 291760 118227 293420 118238
rect 291760 118109 293211 118227
rect 293329 118109 293420 118227
rect 291760 118067 293420 118109
rect 291760 117949 293211 118067
rect 293329 117949 293420 118067
rect 291760 117938 293420 117949
rect -1458 117937 -1158 117938
rect 293120 117937 293420 117938
rect -3758 114638 -3458 114639
rect 295420 114638 295720 114639
rect -4218 114627 240 114638
rect -4218 114509 -3667 114627
rect -3549 114509 240 114627
rect -4218 114467 240 114509
rect -4218 114349 -3667 114467
rect -3549 114349 240 114467
rect -4218 114338 240 114349
rect 291760 114627 296180 114638
rect 291760 114509 295511 114627
rect 295629 114509 296180 114627
rect 291760 114467 296180 114509
rect 291760 114349 295511 114467
rect 295629 114349 296180 114467
rect 291760 114338 296180 114349
rect -3758 114337 -3458 114338
rect 295420 114337 295720 114338
rect -2838 112838 -2538 112839
rect 294500 112838 294800 112839
rect -3298 112827 240 112838
rect -3298 112709 -2747 112827
rect -2629 112709 240 112827
rect -3298 112667 240 112709
rect -3298 112549 -2747 112667
rect -2629 112549 240 112667
rect -3298 112538 240 112549
rect 291760 112827 295260 112838
rect 291760 112709 294591 112827
rect 294709 112709 295260 112827
rect 291760 112667 295260 112709
rect 291760 112549 294591 112667
rect 294709 112549 295260 112667
rect 291760 112538 295260 112549
rect -2838 112537 -2538 112538
rect 294500 112537 294800 112538
rect -1918 111038 -1618 111039
rect 293580 111038 293880 111039
rect -2378 111027 240 111038
rect -2378 110909 -1827 111027
rect -1709 110909 240 111027
rect -2378 110867 240 110909
rect -2378 110749 -1827 110867
rect -1709 110749 240 110867
rect -2378 110738 240 110749
rect 291760 111027 294340 111038
rect 291760 110909 293671 111027
rect 293789 110909 294340 111027
rect 291760 110867 294340 110909
rect 291760 110749 293671 110867
rect 293789 110749 294340 110867
rect 291760 110738 294340 110749
rect -1918 110737 -1618 110738
rect 293580 110737 293880 110738
rect -998 109238 -698 109239
rect 292660 109238 292960 109239
rect -1458 109227 240 109238
rect -1458 109109 -907 109227
rect -789 109109 240 109227
rect -1458 109067 240 109109
rect -1458 108949 -907 109067
rect -789 108949 240 109067
rect -1458 108938 240 108949
rect 291760 109227 293420 109238
rect 291760 109109 292751 109227
rect 292869 109109 293420 109227
rect 291760 109067 293420 109109
rect 291760 108949 292751 109067
rect 292869 108949 293420 109067
rect 291760 108938 293420 108949
rect -998 108937 -698 108938
rect 292660 108937 292960 108938
rect -4218 105638 -3918 105639
rect 295880 105638 296180 105639
rect -4218 105627 240 105638
rect -4218 105509 -4127 105627
rect -4009 105509 240 105627
rect -4218 105467 240 105509
rect -4218 105349 -4127 105467
rect -4009 105349 240 105467
rect -4218 105338 240 105349
rect 291760 105627 296180 105638
rect 291760 105509 295971 105627
rect 296089 105509 296180 105627
rect 291760 105467 296180 105509
rect 291760 105349 295971 105467
rect 296089 105349 296180 105467
rect 291760 105338 296180 105349
rect -4218 105337 -3918 105338
rect 295880 105337 296180 105338
rect -3298 103838 -2998 103839
rect 294960 103838 295260 103839
rect -3298 103827 240 103838
rect -3298 103709 -3207 103827
rect -3089 103709 240 103827
rect -3298 103667 240 103709
rect -3298 103549 -3207 103667
rect -3089 103549 240 103667
rect -3298 103538 240 103549
rect 291760 103827 295260 103838
rect 291760 103709 295051 103827
rect 295169 103709 295260 103827
rect 291760 103667 295260 103709
rect 291760 103549 295051 103667
rect 295169 103549 295260 103667
rect 291760 103538 295260 103549
rect -3298 103537 -2998 103538
rect 294960 103537 295260 103538
rect -2378 102038 -2078 102039
rect 294040 102038 294340 102039
rect -2378 102027 240 102038
rect -2378 101909 -2287 102027
rect -2169 101909 240 102027
rect -2378 101867 240 101909
rect -2378 101749 -2287 101867
rect -2169 101749 240 101867
rect -2378 101738 240 101749
rect 291760 102027 294340 102038
rect 291760 101909 294131 102027
rect 294249 101909 294340 102027
rect 291760 101867 294340 101909
rect 291760 101749 294131 101867
rect 294249 101749 294340 101867
rect 291760 101738 294340 101749
rect -2378 101737 -2078 101738
rect 294040 101737 294340 101738
rect -1458 100238 -1158 100239
rect 293120 100238 293420 100239
rect -1458 100227 240 100238
rect -1458 100109 -1367 100227
rect -1249 100109 240 100227
rect -1458 100067 240 100109
rect -1458 99949 -1367 100067
rect -1249 99949 240 100067
rect -1458 99938 240 99949
rect 291760 100227 293420 100238
rect 291760 100109 293211 100227
rect 293329 100109 293420 100227
rect 291760 100067 293420 100109
rect 291760 99949 293211 100067
rect 293329 99949 293420 100067
rect 291760 99938 293420 99949
rect -1458 99937 -1158 99938
rect 293120 99937 293420 99938
rect -3758 96638 -3458 96639
rect 295420 96638 295720 96639
rect -4218 96627 240 96638
rect -4218 96509 -3667 96627
rect -3549 96509 240 96627
rect -4218 96467 240 96509
rect -4218 96349 -3667 96467
rect -3549 96349 240 96467
rect -4218 96338 240 96349
rect 291760 96627 296180 96638
rect 291760 96509 295511 96627
rect 295629 96509 296180 96627
rect 291760 96467 296180 96509
rect 291760 96349 295511 96467
rect 295629 96349 296180 96467
rect 291760 96338 296180 96349
rect -3758 96337 -3458 96338
rect 295420 96337 295720 96338
rect -2838 94838 -2538 94839
rect 294500 94838 294800 94839
rect -3298 94827 240 94838
rect -3298 94709 -2747 94827
rect -2629 94709 240 94827
rect -3298 94667 240 94709
rect -3298 94549 -2747 94667
rect -2629 94549 240 94667
rect -3298 94538 240 94549
rect 291760 94827 295260 94838
rect 291760 94709 294591 94827
rect 294709 94709 295260 94827
rect 291760 94667 295260 94709
rect 291760 94549 294591 94667
rect 294709 94549 295260 94667
rect 291760 94538 295260 94549
rect -2838 94537 -2538 94538
rect 294500 94537 294800 94538
rect -1918 93038 -1618 93039
rect 293580 93038 293880 93039
rect -2378 93027 240 93038
rect -2378 92909 -1827 93027
rect -1709 92909 240 93027
rect -2378 92867 240 92909
rect -2378 92749 -1827 92867
rect -1709 92749 240 92867
rect -2378 92738 240 92749
rect 291760 93027 294340 93038
rect 291760 92909 293671 93027
rect 293789 92909 294340 93027
rect 291760 92867 294340 92909
rect 291760 92749 293671 92867
rect 293789 92749 294340 92867
rect 291760 92738 294340 92749
rect -1918 92737 -1618 92738
rect 293580 92737 293880 92738
rect -998 91238 -698 91239
rect 292660 91238 292960 91239
rect -1458 91227 240 91238
rect -1458 91109 -907 91227
rect -789 91109 240 91227
rect -1458 91067 240 91109
rect -1458 90949 -907 91067
rect -789 90949 240 91067
rect -1458 90938 240 90949
rect 291760 91227 293420 91238
rect 291760 91109 292751 91227
rect 292869 91109 293420 91227
rect 291760 91067 293420 91109
rect 291760 90949 292751 91067
rect 292869 90949 293420 91067
rect 291760 90938 293420 90949
rect -998 90937 -698 90938
rect 292660 90937 292960 90938
rect -4218 87638 -3918 87639
rect 295880 87638 296180 87639
rect -4218 87627 240 87638
rect -4218 87509 -4127 87627
rect -4009 87509 240 87627
rect -4218 87467 240 87509
rect -4218 87349 -4127 87467
rect -4009 87349 240 87467
rect -4218 87338 240 87349
rect 291760 87627 296180 87638
rect 291760 87509 295971 87627
rect 296089 87509 296180 87627
rect 291760 87467 296180 87509
rect 291760 87349 295971 87467
rect 296089 87349 296180 87467
rect 291760 87338 296180 87349
rect -4218 87337 -3918 87338
rect 295880 87337 296180 87338
rect -3298 85838 -2998 85839
rect 294960 85838 295260 85839
rect -3298 85827 240 85838
rect -3298 85709 -3207 85827
rect -3089 85709 240 85827
rect -3298 85667 240 85709
rect -3298 85549 -3207 85667
rect -3089 85549 240 85667
rect -3298 85538 240 85549
rect 291760 85827 295260 85838
rect 291760 85709 295051 85827
rect 295169 85709 295260 85827
rect 291760 85667 295260 85709
rect 291760 85549 295051 85667
rect 295169 85549 295260 85667
rect 291760 85538 295260 85549
rect -3298 85537 -2998 85538
rect 294960 85537 295260 85538
rect -2378 84038 -2078 84039
rect 294040 84038 294340 84039
rect -2378 84027 240 84038
rect -2378 83909 -2287 84027
rect -2169 83909 240 84027
rect -2378 83867 240 83909
rect -2378 83749 -2287 83867
rect -2169 83749 240 83867
rect -2378 83738 240 83749
rect 291760 84027 294340 84038
rect 291760 83909 294131 84027
rect 294249 83909 294340 84027
rect 291760 83867 294340 83909
rect 291760 83749 294131 83867
rect 294249 83749 294340 83867
rect 291760 83738 294340 83749
rect -2378 83737 -2078 83738
rect 294040 83737 294340 83738
rect -1458 82238 -1158 82239
rect 293120 82238 293420 82239
rect -1458 82227 240 82238
rect -1458 82109 -1367 82227
rect -1249 82109 240 82227
rect -1458 82067 240 82109
rect -1458 81949 -1367 82067
rect -1249 81949 240 82067
rect -1458 81938 240 81949
rect 291760 82227 293420 82238
rect 291760 82109 293211 82227
rect 293329 82109 293420 82227
rect 291760 82067 293420 82109
rect 291760 81949 293211 82067
rect 293329 81949 293420 82067
rect 291760 81938 293420 81949
rect -1458 81937 -1158 81938
rect 293120 81937 293420 81938
rect -3758 78638 -3458 78639
rect 295420 78638 295720 78639
rect -4218 78627 240 78638
rect -4218 78509 -3667 78627
rect -3549 78509 240 78627
rect -4218 78467 240 78509
rect -4218 78349 -3667 78467
rect -3549 78349 240 78467
rect -4218 78338 240 78349
rect 291760 78627 296180 78638
rect 291760 78509 295511 78627
rect 295629 78509 296180 78627
rect 291760 78467 296180 78509
rect 291760 78349 295511 78467
rect 295629 78349 296180 78467
rect 291760 78338 296180 78349
rect -3758 78337 -3458 78338
rect 295420 78337 295720 78338
rect -2838 76838 -2538 76839
rect 294500 76838 294800 76839
rect -3298 76827 240 76838
rect -3298 76709 -2747 76827
rect -2629 76709 240 76827
rect -3298 76667 240 76709
rect -3298 76549 -2747 76667
rect -2629 76549 240 76667
rect -3298 76538 240 76549
rect 291760 76827 295260 76838
rect 291760 76709 294591 76827
rect 294709 76709 295260 76827
rect 291760 76667 295260 76709
rect 291760 76549 294591 76667
rect 294709 76549 295260 76667
rect 291760 76538 295260 76549
rect -2838 76537 -2538 76538
rect 294500 76537 294800 76538
rect -1918 75038 -1618 75039
rect 293580 75038 293880 75039
rect -2378 75027 240 75038
rect -2378 74909 -1827 75027
rect -1709 74909 240 75027
rect -2378 74867 240 74909
rect -2378 74749 -1827 74867
rect -1709 74749 240 74867
rect -2378 74738 240 74749
rect 291760 75027 294340 75038
rect 291760 74909 293671 75027
rect 293789 74909 294340 75027
rect 291760 74867 294340 74909
rect 291760 74749 293671 74867
rect 293789 74749 294340 74867
rect 291760 74738 294340 74749
rect -1918 74737 -1618 74738
rect 293580 74737 293880 74738
rect -998 73238 -698 73239
rect 292660 73238 292960 73239
rect -1458 73227 240 73238
rect -1458 73109 -907 73227
rect -789 73109 240 73227
rect -1458 73067 240 73109
rect -1458 72949 -907 73067
rect -789 72949 240 73067
rect -1458 72938 240 72949
rect 291760 73227 293420 73238
rect 291760 73109 292751 73227
rect 292869 73109 293420 73227
rect 291760 73067 293420 73109
rect 291760 72949 292751 73067
rect 292869 72949 293420 73067
rect 291760 72938 293420 72949
rect -998 72937 -698 72938
rect 292660 72937 292960 72938
rect -4218 69638 -3918 69639
rect 295880 69638 296180 69639
rect -4218 69627 240 69638
rect -4218 69509 -4127 69627
rect -4009 69509 240 69627
rect -4218 69467 240 69509
rect -4218 69349 -4127 69467
rect -4009 69349 240 69467
rect -4218 69338 240 69349
rect 291760 69627 296180 69638
rect 291760 69509 295971 69627
rect 296089 69509 296180 69627
rect 291760 69467 296180 69509
rect 291760 69349 295971 69467
rect 296089 69349 296180 69467
rect 291760 69338 296180 69349
rect -4218 69337 -3918 69338
rect 295880 69337 296180 69338
rect -3298 67838 -2998 67839
rect 294960 67838 295260 67839
rect -3298 67827 240 67838
rect -3298 67709 -3207 67827
rect -3089 67709 240 67827
rect -3298 67667 240 67709
rect -3298 67549 -3207 67667
rect -3089 67549 240 67667
rect -3298 67538 240 67549
rect 291760 67827 295260 67838
rect 291760 67709 295051 67827
rect 295169 67709 295260 67827
rect 291760 67667 295260 67709
rect 291760 67549 295051 67667
rect 295169 67549 295260 67667
rect 291760 67538 295260 67549
rect -3298 67537 -2998 67538
rect 294960 67537 295260 67538
rect -2378 66038 -2078 66039
rect 294040 66038 294340 66039
rect -2378 66027 240 66038
rect -2378 65909 -2287 66027
rect -2169 65909 240 66027
rect -2378 65867 240 65909
rect -2378 65749 -2287 65867
rect -2169 65749 240 65867
rect -2378 65738 240 65749
rect 291760 66027 294340 66038
rect 291760 65909 294131 66027
rect 294249 65909 294340 66027
rect 291760 65867 294340 65909
rect 291760 65749 294131 65867
rect 294249 65749 294340 65867
rect 291760 65738 294340 65749
rect -2378 65737 -2078 65738
rect 294040 65737 294340 65738
rect -1458 64238 -1158 64239
rect 293120 64238 293420 64239
rect -1458 64227 240 64238
rect -1458 64109 -1367 64227
rect -1249 64109 240 64227
rect -1458 64067 240 64109
rect -1458 63949 -1367 64067
rect -1249 63949 240 64067
rect -1458 63938 240 63949
rect 291760 64227 293420 64238
rect 291760 64109 293211 64227
rect 293329 64109 293420 64227
rect 291760 64067 293420 64109
rect 291760 63949 293211 64067
rect 293329 63949 293420 64067
rect 291760 63938 293420 63949
rect -1458 63937 -1158 63938
rect 293120 63937 293420 63938
rect -3758 60638 -3458 60639
rect 295420 60638 295720 60639
rect -4218 60627 240 60638
rect -4218 60509 -3667 60627
rect -3549 60509 240 60627
rect -4218 60467 240 60509
rect -4218 60349 -3667 60467
rect -3549 60349 240 60467
rect -4218 60338 240 60349
rect 291760 60627 296180 60638
rect 291760 60509 295511 60627
rect 295629 60509 296180 60627
rect 291760 60467 296180 60509
rect 291760 60349 295511 60467
rect 295629 60349 296180 60467
rect 291760 60338 296180 60349
rect -3758 60337 -3458 60338
rect 295420 60337 295720 60338
rect -2838 58838 -2538 58839
rect 294500 58838 294800 58839
rect -3298 58827 240 58838
rect -3298 58709 -2747 58827
rect -2629 58709 240 58827
rect -3298 58667 240 58709
rect -3298 58549 -2747 58667
rect -2629 58549 240 58667
rect -3298 58538 240 58549
rect 291760 58827 295260 58838
rect 291760 58709 294591 58827
rect 294709 58709 295260 58827
rect 291760 58667 295260 58709
rect 291760 58549 294591 58667
rect 294709 58549 295260 58667
rect 291760 58538 295260 58549
rect -2838 58537 -2538 58538
rect 294500 58537 294800 58538
rect -1918 57038 -1618 57039
rect 293580 57038 293880 57039
rect -2378 57027 240 57038
rect -2378 56909 -1827 57027
rect -1709 56909 240 57027
rect -2378 56867 240 56909
rect -2378 56749 -1827 56867
rect -1709 56749 240 56867
rect -2378 56738 240 56749
rect 291760 57027 294340 57038
rect 291760 56909 293671 57027
rect 293789 56909 294340 57027
rect 291760 56867 294340 56909
rect 291760 56749 293671 56867
rect 293789 56749 294340 56867
rect 291760 56738 294340 56749
rect -1918 56737 -1618 56738
rect 293580 56737 293880 56738
rect -998 55238 -698 55239
rect 292660 55238 292960 55239
rect -1458 55227 240 55238
rect -1458 55109 -907 55227
rect -789 55109 240 55227
rect -1458 55067 240 55109
rect -1458 54949 -907 55067
rect -789 54949 240 55067
rect -1458 54938 240 54949
rect 291760 55227 293420 55238
rect 291760 55109 292751 55227
rect 292869 55109 293420 55227
rect 291760 55067 293420 55109
rect 291760 54949 292751 55067
rect 292869 54949 293420 55067
rect 291760 54938 293420 54949
rect -998 54937 -698 54938
rect 292660 54937 292960 54938
rect -4218 51638 -3918 51639
rect 295880 51638 296180 51639
rect -4218 51627 240 51638
rect -4218 51509 -4127 51627
rect -4009 51509 240 51627
rect -4218 51467 240 51509
rect -4218 51349 -4127 51467
rect -4009 51349 240 51467
rect -4218 51338 240 51349
rect 291760 51627 296180 51638
rect 291760 51509 295971 51627
rect 296089 51509 296180 51627
rect 291760 51467 296180 51509
rect 291760 51349 295971 51467
rect 296089 51349 296180 51467
rect 291760 51338 296180 51349
rect -4218 51337 -3918 51338
rect 295880 51337 296180 51338
rect -3298 49838 -2998 49839
rect 294960 49838 295260 49839
rect -3298 49827 240 49838
rect -3298 49709 -3207 49827
rect -3089 49709 240 49827
rect -3298 49667 240 49709
rect -3298 49549 -3207 49667
rect -3089 49549 240 49667
rect -3298 49538 240 49549
rect 291760 49827 295260 49838
rect 291760 49709 295051 49827
rect 295169 49709 295260 49827
rect 291760 49667 295260 49709
rect 291760 49549 295051 49667
rect 295169 49549 295260 49667
rect 291760 49538 295260 49549
rect -3298 49537 -2998 49538
rect 294960 49537 295260 49538
rect -2378 48038 -2078 48039
rect 294040 48038 294340 48039
rect -2378 48027 240 48038
rect -2378 47909 -2287 48027
rect -2169 47909 240 48027
rect -2378 47867 240 47909
rect -2378 47749 -2287 47867
rect -2169 47749 240 47867
rect -2378 47738 240 47749
rect 291760 48027 294340 48038
rect 291760 47909 294131 48027
rect 294249 47909 294340 48027
rect 291760 47867 294340 47909
rect 291760 47749 294131 47867
rect 294249 47749 294340 47867
rect 291760 47738 294340 47749
rect -2378 47737 -2078 47738
rect 294040 47737 294340 47738
rect -1458 46238 -1158 46239
rect 293120 46238 293420 46239
rect -1458 46227 240 46238
rect -1458 46109 -1367 46227
rect -1249 46109 240 46227
rect -1458 46067 240 46109
rect -1458 45949 -1367 46067
rect -1249 45949 240 46067
rect -1458 45938 240 45949
rect 291760 46227 293420 46238
rect 291760 46109 293211 46227
rect 293329 46109 293420 46227
rect 291760 46067 293420 46109
rect 291760 45949 293211 46067
rect 293329 45949 293420 46067
rect 291760 45938 293420 45949
rect -1458 45937 -1158 45938
rect 293120 45937 293420 45938
rect -3758 42638 -3458 42639
rect 295420 42638 295720 42639
rect -4218 42627 240 42638
rect -4218 42509 -3667 42627
rect -3549 42509 240 42627
rect -4218 42467 240 42509
rect -4218 42349 -3667 42467
rect -3549 42349 240 42467
rect -4218 42338 240 42349
rect 291760 42627 296180 42638
rect 291760 42509 295511 42627
rect 295629 42509 296180 42627
rect 291760 42467 296180 42509
rect 291760 42349 295511 42467
rect 295629 42349 296180 42467
rect 291760 42338 296180 42349
rect -3758 42337 -3458 42338
rect 295420 42337 295720 42338
rect -2838 40838 -2538 40839
rect 294500 40838 294800 40839
rect -3298 40827 240 40838
rect -3298 40709 -2747 40827
rect -2629 40709 240 40827
rect -3298 40667 240 40709
rect -3298 40549 -2747 40667
rect -2629 40549 240 40667
rect -3298 40538 240 40549
rect 291760 40827 295260 40838
rect 291760 40709 294591 40827
rect 294709 40709 295260 40827
rect 291760 40667 295260 40709
rect 291760 40549 294591 40667
rect 294709 40549 295260 40667
rect 291760 40538 295260 40549
rect -2838 40537 -2538 40538
rect 294500 40537 294800 40538
rect -1918 39038 -1618 39039
rect 293580 39038 293880 39039
rect -2378 39027 240 39038
rect -2378 38909 -1827 39027
rect -1709 38909 240 39027
rect -2378 38867 240 38909
rect -2378 38749 -1827 38867
rect -1709 38749 240 38867
rect -2378 38738 240 38749
rect 291760 39027 294340 39038
rect 291760 38909 293671 39027
rect 293789 38909 294340 39027
rect 291760 38867 294340 38909
rect 291760 38749 293671 38867
rect 293789 38749 294340 38867
rect 291760 38738 294340 38749
rect -1918 38737 -1618 38738
rect 293580 38737 293880 38738
rect -998 37238 -698 37239
rect 292660 37238 292960 37239
rect -1458 37227 240 37238
rect -1458 37109 -907 37227
rect -789 37109 240 37227
rect -1458 37067 240 37109
rect -1458 36949 -907 37067
rect -789 36949 240 37067
rect -1458 36938 240 36949
rect 291760 37227 293420 37238
rect 291760 37109 292751 37227
rect 292869 37109 293420 37227
rect 291760 37067 293420 37109
rect 291760 36949 292751 37067
rect 292869 36949 293420 37067
rect 291760 36938 293420 36949
rect -998 36937 -698 36938
rect 292660 36937 292960 36938
rect -4218 33638 -3918 33639
rect 295880 33638 296180 33639
rect -4218 33627 240 33638
rect -4218 33509 -4127 33627
rect -4009 33509 240 33627
rect -4218 33467 240 33509
rect -4218 33349 -4127 33467
rect -4009 33349 240 33467
rect -4218 33338 240 33349
rect 291760 33627 296180 33638
rect 291760 33509 295971 33627
rect 296089 33509 296180 33627
rect 291760 33467 296180 33509
rect 291760 33349 295971 33467
rect 296089 33349 296180 33467
rect 291760 33338 296180 33349
rect -4218 33337 -3918 33338
rect 295880 33337 296180 33338
rect -3298 31838 -2998 31839
rect 294960 31838 295260 31839
rect -3298 31827 240 31838
rect -3298 31709 -3207 31827
rect -3089 31709 240 31827
rect -3298 31667 240 31709
rect -3298 31549 -3207 31667
rect -3089 31549 240 31667
rect -3298 31538 240 31549
rect 291760 31827 295260 31838
rect 291760 31709 295051 31827
rect 295169 31709 295260 31827
rect 291760 31667 295260 31709
rect 291760 31549 295051 31667
rect 295169 31549 295260 31667
rect 291760 31538 295260 31549
rect -3298 31537 -2998 31538
rect 294960 31537 295260 31538
rect -2378 30038 -2078 30039
rect 294040 30038 294340 30039
rect -2378 30027 240 30038
rect -2378 29909 -2287 30027
rect -2169 29909 240 30027
rect -2378 29867 240 29909
rect -2378 29749 -2287 29867
rect -2169 29749 240 29867
rect -2378 29738 240 29749
rect 291760 30027 294340 30038
rect 291760 29909 294131 30027
rect 294249 29909 294340 30027
rect 291760 29867 294340 29909
rect 291760 29749 294131 29867
rect 294249 29749 294340 29867
rect 291760 29738 294340 29749
rect -2378 29737 -2078 29738
rect 294040 29737 294340 29738
rect -1458 28238 -1158 28239
rect 293120 28238 293420 28239
rect -1458 28227 240 28238
rect -1458 28109 -1367 28227
rect -1249 28109 240 28227
rect -1458 28067 240 28109
rect -1458 27949 -1367 28067
rect -1249 27949 240 28067
rect -1458 27938 240 27949
rect 291760 28227 293420 28238
rect 291760 28109 293211 28227
rect 293329 28109 293420 28227
rect 291760 28067 293420 28109
rect 291760 27949 293211 28067
rect 293329 27949 293420 28067
rect 291760 27938 293420 27949
rect -1458 27937 -1158 27938
rect 293120 27937 293420 27938
rect -3758 24638 -3458 24639
rect 295420 24638 295720 24639
rect -4218 24627 240 24638
rect -4218 24509 -3667 24627
rect -3549 24509 240 24627
rect -4218 24467 240 24509
rect -4218 24349 -3667 24467
rect -3549 24349 240 24467
rect -4218 24338 240 24349
rect 291760 24627 296180 24638
rect 291760 24509 295511 24627
rect 295629 24509 296180 24627
rect 291760 24467 296180 24509
rect 291760 24349 295511 24467
rect 295629 24349 296180 24467
rect 291760 24338 296180 24349
rect -3758 24337 -3458 24338
rect 295420 24337 295720 24338
rect -2838 22838 -2538 22839
rect 294500 22838 294800 22839
rect -3298 22827 240 22838
rect -3298 22709 -2747 22827
rect -2629 22709 240 22827
rect -3298 22667 240 22709
rect -3298 22549 -2747 22667
rect -2629 22549 240 22667
rect -3298 22538 240 22549
rect 291760 22827 295260 22838
rect 291760 22709 294591 22827
rect 294709 22709 295260 22827
rect 291760 22667 295260 22709
rect 291760 22549 294591 22667
rect 294709 22549 295260 22667
rect 291760 22538 295260 22549
rect -2838 22537 -2538 22538
rect 294500 22537 294800 22538
rect -1918 21038 -1618 21039
rect 293580 21038 293880 21039
rect -2378 21027 240 21038
rect -2378 20909 -1827 21027
rect -1709 20909 240 21027
rect -2378 20867 240 20909
rect -2378 20749 -1827 20867
rect -1709 20749 240 20867
rect -2378 20738 240 20749
rect 291760 21027 294340 21038
rect 291760 20909 293671 21027
rect 293789 20909 294340 21027
rect 291760 20867 294340 20909
rect 291760 20749 293671 20867
rect 293789 20749 294340 20867
rect 291760 20738 294340 20749
rect -1918 20737 -1618 20738
rect 293580 20737 293880 20738
rect -998 19238 -698 19239
rect 292660 19238 292960 19239
rect -1458 19227 240 19238
rect -1458 19109 -907 19227
rect -789 19109 240 19227
rect -1458 19067 240 19109
rect -1458 18949 -907 19067
rect -789 18949 240 19067
rect -1458 18938 240 18949
rect 291760 19227 293420 19238
rect 291760 19109 292751 19227
rect 292869 19109 293420 19227
rect 291760 19067 293420 19109
rect 291760 18949 292751 19067
rect 292869 18949 293420 19067
rect 291760 18938 293420 18949
rect -998 18937 -698 18938
rect 292660 18937 292960 18938
rect -4218 15638 -3918 15639
rect 295880 15638 296180 15639
rect -4218 15627 240 15638
rect -4218 15509 -4127 15627
rect -4009 15509 240 15627
rect -4218 15467 240 15509
rect -4218 15349 -4127 15467
rect -4009 15349 240 15467
rect -4218 15338 240 15349
rect 291760 15627 296180 15638
rect 291760 15509 295971 15627
rect 296089 15509 296180 15627
rect 291760 15467 296180 15509
rect 291760 15349 295971 15467
rect 296089 15349 296180 15467
rect 291760 15338 296180 15349
rect -4218 15337 -3918 15338
rect 295880 15337 296180 15338
rect -3298 13838 -2998 13839
rect 294960 13838 295260 13839
rect -3298 13827 240 13838
rect -3298 13709 -3207 13827
rect -3089 13709 240 13827
rect -3298 13667 240 13709
rect -3298 13549 -3207 13667
rect -3089 13549 240 13667
rect -3298 13538 240 13549
rect 291760 13827 295260 13838
rect 291760 13709 295051 13827
rect 295169 13709 295260 13827
rect 291760 13667 295260 13709
rect 291760 13549 295051 13667
rect 295169 13549 295260 13667
rect 291760 13538 295260 13549
rect -3298 13537 -2998 13538
rect 294960 13537 295260 13538
rect -2378 12038 -2078 12039
rect 294040 12038 294340 12039
rect -2378 12027 240 12038
rect -2378 11909 -2287 12027
rect -2169 11909 240 12027
rect -2378 11867 240 11909
rect -2378 11749 -2287 11867
rect -2169 11749 240 11867
rect -2378 11738 240 11749
rect 291760 12027 294340 12038
rect 291760 11909 294131 12027
rect 294249 11909 294340 12027
rect 291760 11867 294340 11909
rect 291760 11749 294131 11867
rect 294249 11749 294340 11867
rect 291760 11738 294340 11749
rect -2378 11737 -2078 11738
rect 294040 11737 294340 11738
rect -1458 10238 -1158 10239
rect 293120 10238 293420 10239
rect -1458 10227 240 10238
rect -1458 10109 -1367 10227
rect -1249 10109 240 10227
rect -1458 10067 240 10109
rect -1458 9949 -1367 10067
rect -1249 9949 240 10067
rect -1458 9938 240 9949
rect 291760 10227 293420 10238
rect 291760 10109 293211 10227
rect 293329 10109 293420 10227
rect 291760 10067 293420 10109
rect 291760 9949 293211 10067
rect 293329 9949 293420 10067
rect 291760 9938 293420 9949
rect -1458 9937 -1158 9938
rect 293120 9937 293420 9938
rect -3758 6638 -3458 6639
rect 295420 6638 295720 6639
rect -4218 6627 240 6638
rect -4218 6509 -3667 6627
rect -3549 6509 240 6627
rect -4218 6467 240 6509
rect -4218 6349 -3667 6467
rect -3549 6349 240 6467
rect -4218 6338 240 6349
rect 291760 6627 296180 6638
rect 291760 6509 295511 6627
rect 295629 6509 296180 6627
rect 291760 6467 296180 6509
rect 291760 6349 295511 6467
rect 295629 6349 296180 6467
rect 291760 6338 296180 6349
rect -3758 6337 -3458 6338
rect 295420 6337 295720 6338
rect -2838 4838 -2538 4839
rect 294500 4838 294800 4839
rect -3298 4827 240 4838
rect -3298 4709 -2747 4827
rect -2629 4709 240 4827
rect -3298 4667 240 4709
rect -3298 4549 -2747 4667
rect -2629 4549 240 4667
rect -3298 4538 240 4549
rect 291760 4827 295260 4838
rect 291760 4709 294591 4827
rect 294709 4709 295260 4827
rect 291760 4667 295260 4709
rect 291760 4549 294591 4667
rect 294709 4549 295260 4667
rect 291760 4538 295260 4549
rect -2838 4537 -2538 4538
rect 294500 4537 294800 4538
rect -1918 3038 -1618 3039
rect 293580 3038 293880 3039
rect -2378 3027 240 3038
rect -2378 2909 -1827 3027
rect -1709 2909 240 3027
rect -2378 2867 240 2909
rect -2378 2749 -1827 2867
rect -1709 2749 240 2867
rect -2378 2738 240 2749
rect 291760 3027 294340 3038
rect 291760 2909 293671 3027
rect 293789 2909 294340 3027
rect 291760 2867 294340 2909
rect 291760 2749 293671 2867
rect 293789 2749 294340 2867
rect 291760 2738 294340 2749
rect -1918 2737 -1618 2738
rect 293580 2737 293880 2738
rect -998 1238 -698 1239
rect 292660 1238 292960 1239
rect -1458 1227 240 1238
rect -1458 1109 -907 1227
rect -789 1109 240 1227
rect -1458 1067 240 1109
rect -1458 949 -907 1067
rect -789 949 240 1067
rect -1458 938 240 949
rect 291760 1227 293420 1238
rect 291760 1109 292751 1227
rect 292869 1109 293420 1227
rect 291760 1067 293420 1109
rect 291760 949 292751 1067
rect 292869 949 293420 1067
rect 291760 938 293420 949
rect -998 937 -698 938
rect 292660 937 292960 938
rect -998 -162 -698 -161
rect 402 -162 702 -161
rect 18402 -162 18702 -161
rect 36402 -162 36702 -161
rect 54402 -162 54702 -161
rect 72402 -162 72702 -161
rect 90402 -162 90702 -161
rect 108402 -162 108702 -161
rect 126402 -162 126702 -161
rect 144402 -162 144702 -161
rect 162402 -162 162702 -161
rect 180402 -162 180702 -161
rect 198402 -162 198702 -161
rect 216402 -162 216702 -161
rect 234402 -162 234702 -161
rect 252402 -162 252702 -161
rect 270402 -162 270702 -161
rect 288402 -162 288702 -161
rect 292660 -162 292960 -161
rect -998 -173 292960 -162
rect -998 -291 -907 -173
rect -789 -291 493 -173
rect 611 -291 18493 -173
rect 18611 -291 36493 -173
rect 36611 -291 54493 -173
rect 54611 -291 72493 -173
rect 72611 -291 90493 -173
rect 90611 -291 108493 -173
rect 108611 -291 126493 -173
rect 126611 -291 144493 -173
rect 144611 -291 162493 -173
rect 162611 -291 180493 -173
rect 180611 -291 198493 -173
rect 198611 -291 216493 -173
rect 216611 -291 234493 -173
rect 234611 -291 252493 -173
rect 252611 -291 270493 -173
rect 270611 -291 288493 -173
rect 288611 -291 292751 -173
rect 292869 -291 292960 -173
rect -998 -333 292960 -291
rect -998 -451 -907 -333
rect -789 -451 493 -333
rect 611 -451 18493 -333
rect 18611 -451 36493 -333
rect 36611 -451 54493 -333
rect 54611 -451 72493 -333
rect 72611 -451 90493 -333
rect 90611 -451 108493 -333
rect 108611 -451 126493 -333
rect 126611 -451 144493 -333
rect 144611 -451 162493 -333
rect 162611 -451 180493 -333
rect 180611 -451 198493 -333
rect 198611 -451 216493 -333
rect 216611 -451 234493 -333
rect 234611 -451 252493 -333
rect 252611 -451 270493 -333
rect 270611 -451 288493 -333
rect 288611 -451 292751 -333
rect 292869 -451 292960 -333
rect -998 -462 292960 -451
rect -998 -463 -698 -462
rect 402 -463 702 -462
rect 18402 -463 18702 -462
rect 36402 -463 36702 -462
rect 54402 -463 54702 -462
rect 72402 -463 72702 -462
rect 90402 -463 90702 -462
rect 108402 -463 108702 -462
rect 126402 -463 126702 -462
rect 144402 -463 144702 -462
rect 162402 -463 162702 -462
rect 180402 -463 180702 -462
rect 198402 -463 198702 -462
rect 216402 -463 216702 -462
rect 234402 -463 234702 -462
rect 252402 -463 252702 -462
rect 270402 -463 270702 -462
rect 288402 -463 288702 -462
rect 292660 -463 292960 -462
rect -1458 -622 -1158 -621
rect 9402 -622 9702 -621
rect 27402 -622 27702 -621
rect 45402 -622 45702 -621
rect 63402 -622 63702 -621
rect 81402 -622 81702 -621
rect 99402 -622 99702 -621
rect 117402 -622 117702 -621
rect 135402 -622 135702 -621
rect 153402 -622 153702 -621
rect 171402 -622 171702 -621
rect 189402 -622 189702 -621
rect 207402 -622 207702 -621
rect 225402 -622 225702 -621
rect 243402 -622 243702 -621
rect 261402 -622 261702 -621
rect 279402 -622 279702 -621
rect 293120 -622 293420 -621
rect -1458 -633 293420 -622
rect -1458 -751 -1367 -633
rect -1249 -751 9493 -633
rect 9611 -751 27493 -633
rect 27611 -751 45493 -633
rect 45611 -751 63493 -633
rect 63611 -751 81493 -633
rect 81611 -751 99493 -633
rect 99611 -751 117493 -633
rect 117611 -751 135493 -633
rect 135611 -751 153493 -633
rect 153611 -751 171493 -633
rect 171611 -751 189493 -633
rect 189611 -751 207493 -633
rect 207611 -751 225493 -633
rect 225611 -751 243493 -633
rect 243611 -751 261493 -633
rect 261611 -751 279493 -633
rect 279611 -751 293211 -633
rect 293329 -751 293420 -633
rect -1458 -793 293420 -751
rect -1458 -911 -1367 -793
rect -1249 -911 9493 -793
rect 9611 -911 27493 -793
rect 27611 -911 45493 -793
rect 45611 -911 63493 -793
rect 63611 -911 81493 -793
rect 81611 -911 99493 -793
rect 99611 -911 117493 -793
rect 117611 -911 135493 -793
rect 135611 -911 153493 -793
rect 153611 -911 171493 -793
rect 171611 -911 189493 -793
rect 189611 -911 207493 -793
rect 207611 -911 225493 -793
rect 225611 -911 243493 -793
rect 243611 -911 261493 -793
rect 261611 -911 279493 -793
rect 279611 -911 293211 -793
rect 293329 -911 293420 -793
rect -1458 -922 293420 -911
rect -1458 -923 -1158 -922
rect 9402 -923 9702 -922
rect 27402 -923 27702 -922
rect 45402 -923 45702 -922
rect 63402 -923 63702 -922
rect 81402 -923 81702 -922
rect 99402 -923 99702 -922
rect 117402 -923 117702 -922
rect 135402 -923 135702 -922
rect 153402 -923 153702 -922
rect 171402 -923 171702 -922
rect 189402 -923 189702 -922
rect 207402 -923 207702 -922
rect 225402 -923 225702 -922
rect 243402 -923 243702 -922
rect 261402 -923 261702 -922
rect 279402 -923 279702 -922
rect 293120 -923 293420 -922
rect -1918 -1082 -1618 -1081
rect 2202 -1082 2502 -1081
rect 20202 -1082 20502 -1081
rect 38202 -1082 38502 -1081
rect 56202 -1082 56502 -1081
rect 74202 -1082 74502 -1081
rect 92202 -1082 92502 -1081
rect 110202 -1082 110502 -1081
rect 128202 -1082 128502 -1081
rect 146202 -1082 146502 -1081
rect 164202 -1082 164502 -1081
rect 182202 -1082 182502 -1081
rect 200202 -1082 200502 -1081
rect 218202 -1082 218502 -1081
rect 236202 -1082 236502 -1081
rect 254202 -1082 254502 -1081
rect 272202 -1082 272502 -1081
rect 290202 -1082 290502 -1081
rect 293580 -1082 293880 -1081
rect -1918 -1093 293880 -1082
rect -1918 -1211 -1827 -1093
rect -1709 -1211 2293 -1093
rect 2411 -1211 20293 -1093
rect 20411 -1211 38293 -1093
rect 38411 -1211 56293 -1093
rect 56411 -1211 74293 -1093
rect 74411 -1211 92293 -1093
rect 92411 -1211 110293 -1093
rect 110411 -1211 128293 -1093
rect 128411 -1211 146293 -1093
rect 146411 -1211 164293 -1093
rect 164411 -1211 182293 -1093
rect 182411 -1211 200293 -1093
rect 200411 -1211 218293 -1093
rect 218411 -1211 236293 -1093
rect 236411 -1211 254293 -1093
rect 254411 -1211 272293 -1093
rect 272411 -1211 290293 -1093
rect 290411 -1211 293671 -1093
rect 293789 -1211 293880 -1093
rect -1918 -1253 293880 -1211
rect -1918 -1371 -1827 -1253
rect -1709 -1371 2293 -1253
rect 2411 -1371 20293 -1253
rect 20411 -1371 38293 -1253
rect 38411 -1371 56293 -1253
rect 56411 -1371 74293 -1253
rect 74411 -1371 92293 -1253
rect 92411 -1371 110293 -1253
rect 110411 -1371 128293 -1253
rect 128411 -1371 146293 -1253
rect 146411 -1371 164293 -1253
rect 164411 -1371 182293 -1253
rect 182411 -1371 200293 -1253
rect 200411 -1371 218293 -1253
rect 218411 -1371 236293 -1253
rect 236411 -1371 254293 -1253
rect 254411 -1371 272293 -1253
rect 272411 -1371 290293 -1253
rect 290411 -1371 293671 -1253
rect 293789 -1371 293880 -1253
rect -1918 -1382 293880 -1371
rect -1918 -1383 -1618 -1382
rect 2202 -1383 2502 -1382
rect 20202 -1383 20502 -1382
rect 38202 -1383 38502 -1382
rect 56202 -1383 56502 -1382
rect 74202 -1383 74502 -1382
rect 92202 -1383 92502 -1382
rect 110202 -1383 110502 -1382
rect 128202 -1383 128502 -1382
rect 146202 -1383 146502 -1382
rect 164202 -1383 164502 -1382
rect 182202 -1383 182502 -1382
rect 200202 -1383 200502 -1382
rect 218202 -1383 218502 -1382
rect 236202 -1383 236502 -1382
rect 254202 -1383 254502 -1382
rect 272202 -1383 272502 -1382
rect 290202 -1383 290502 -1382
rect 293580 -1383 293880 -1382
rect -2378 -1542 -2078 -1541
rect 11202 -1542 11502 -1541
rect 29202 -1542 29502 -1541
rect 47202 -1542 47502 -1541
rect 65202 -1542 65502 -1541
rect 83202 -1542 83502 -1541
rect 101202 -1542 101502 -1541
rect 119202 -1542 119502 -1541
rect 137202 -1542 137502 -1541
rect 155202 -1542 155502 -1541
rect 173202 -1542 173502 -1541
rect 191202 -1542 191502 -1541
rect 209202 -1542 209502 -1541
rect 227202 -1542 227502 -1541
rect 245202 -1542 245502 -1541
rect 263202 -1542 263502 -1541
rect 281202 -1542 281502 -1541
rect 294040 -1542 294340 -1541
rect -2378 -1553 294340 -1542
rect -2378 -1671 -2287 -1553
rect -2169 -1671 11293 -1553
rect 11411 -1671 29293 -1553
rect 29411 -1671 47293 -1553
rect 47411 -1671 65293 -1553
rect 65411 -1671 83293 -1553
rect 83411 -1671 101293 -1553
rect 101411 -1671 119293 -1553
rect 119411 -1671 137293 -1553
rect 137411 -1671 155293 -1553
rect 155411 -1671 173293 -1553
rect 173411 -1671 191293 -1553
rect 191411 -1671 209293 -1553
rect 209411 -1671 227293 -1553
rect 227411 -1671 245293 -1553
rect 245411 -1671 263293 -1553
rect 263411 -1671 281293 -1553
rect 281411 -1671 294131 -1553
rect 294249 -1671 294340 -1553
rect -2378 -1713 294340 -1671
rect -2378 -1831 -2287 -1713
rect -2169 -1831 11293 -1713
rect 11411 -1831 29293 -1713
rect 29411 -1831 47293 -1713
rect 47411 -1831 65293 -1713
rect 65411 -1831 83293 -1713
rect 83411 -1831 101293 -1713
rect 101411 -1831 119293 -1713
rect 119411 -1831 137293 -1713
rect 137411 -1831 155293 -1713
rect 155411 -1831 173293 -1713
rect 173411 -1831 191293 -1713
rect 191411 -1831 209293 -1713
rect 209411 -1831 227293 -1713
rect 227411 -1831 245293 -1713
rect 245411 -1831 263293 -1713
rect 263411 -1831 281293 -1713
rect 281411 -1831 294131 -1713
rect 294249 -1831 294340 -1713
rect -2378 -1842 294340 -1831
rect -2378 -1843 -2078 -1842
rect 11202 -1843 11502 -1842
rect 29202 -1843 29502 -1842
rect 47202 -1843 47502 -1842
rect 65202 -1843 65502 -1842
rect 83202 -1843 83502 -1842
rect 101202 -1843 101502 -1842
rect 119202 -1843 119502 -1842
rect 137202 -1843 137502 -1842
rect 155202 -1843 155502 -1842
rect 173202 -1843 173502 -1842
rect 191202 -1843 191502 -1842
rect 209202 -1843 209502 -1842
rect 227202 -1843 227502 -1842
rect 245202 -1843 245502 -1842
rect 263202 -1843 263502 -1842
rect 281202 -1843 281502 -1842
rect 294040 -1843 294340 -1842
rect -2838 -2002 -2538 -2001
rect 4002 -2002 4302 -2001
rect 22002 -2002 22302 -2001
rect 40002 -2002 40302 -2001
rect 58002 -2002 58302 -2001
rect 76002 -2002 76302 -2001
rect 94002 -2002 94302 -2001
rect 112002 -2002 112302 -2001
rect 130002 -2002 130302 -2001
rect 148002 -2002 148302 -2001
rect 166002 -2002 166302 -2001
rect 184002 -2002 184302 -2001
rect 202002 -2002 202302 -2001
rect 220002 -2002 220302 -2001
rect 238002 -2002 238302 -2001
rect 256002 -2002 256302 -2001
rect 274002 -2002 274302 -2001
rect 294500 -2002 294800 -2001
rect -2838 -2013 294800 -2002
rect -2838 -2131 -2747 -2013
rect -2629 -2131 4093 -2013
rect 4211 -2131 22093 -2013
rect 22211 -2131 40093 -2013
rect 40211 -2131 58093 -2013
rect 58211 -2131 76093 -2013
rect 76211 -2131 94093 -2013
rect 94211 -2131 112093 -2013
rect 112211 -2131 130093 -2013
rect 130211 -2131 148093 -2013
rect 148211 -2131 166093 -2013
rect 166211 -2131 184093 -2013
rect 184211 -2131 202093 -2013
rect 202211 -2131 220093 -2013
rect 220211 -2131 238093 -2013
rect 238211 -2131 256093 -2013
rect 256211 -2131 274093 -2013
rect 274211 -2131 294591 -2013
rect 294709 -2131 294800 -2013
rect -2838 -2173 294800 -2131
rect -2838 -2291 -2747 -2173
rect -2629 -2291 4093 -2173
rect 4211 -2291 22093 -2173
rect 22211 -2291 40093 -2173
rect 40211 -2291 58093 -2173
rect 58211 -2291 76093 -2173
rect 76211 -2291 94093 -2173
rect 94211 -2291 112093 -2173
rect 112211 -2291 130093 -2173
rect 130211 -2291 148093 -2173
rect 148211 -2291 166093 -2173
rect 166211 -2291 184093 -2173
rect 184211 -2291 202093 -2173
rect 202211 -2291 220093 -2173
rect 220211 -2291 238093 -2173
rect 238211 -2291 256093 -2173
rect 256211 -2291 274093 -2173
rect 274211 -2291 294591 -2173
rect 294709 -2291 294800 -2173
rect -2838 -2302 294800 -2291
rect -2838 -2303 -2538 -2302
rect 4002 -2303 4302 -2302
rect 22002 -2303 22302 -2302
rect 40002 -2303 40302 -2302
rect 58002 -2303 58302 -2302
rect 76002 -2303 76302 -2302
rect 94002 -2303 94302 -2302
rect 112002 -2303 112302 -2302
rect 130002 -2303 130302 -2302
rect 148002 -2303 148302 -2302
rect 166002 -2303 166302 -2302
rect 184002 -2303 184302 -2302
rect 202002 -2303 202302 -2302
rect 220002 -2303 220302 -2302
rect 238002 -2303 238302 -2302
rect 256002 -2303 256302 -2302
rect 274002 -2303 274302 -2302
rect 294500 -2303 294800 -2302
rect -3298 -2462 -2998 -2461
rect 13002 -2462 13302 -2461
rect 31002 -2462 31302 -2461
rect 49002 -2462 49302 -2461
rect 67002 -2462 67302 -2461
rect 85002 -2462 85302 -2461
rect 103002 -2462 103302 -2461
rect 121002 -2462 121302 -2461
rect 139002 -2462 139302 -2461
rect 157002 -2462 157302 -2461
rect 175002 -2462 175302 -2461
rect 193002 -2462 193302 -2461
rect 211002 -2462 211302 -2461
rect 229002 -2462 229302 -2461
rect 247002 -2462 247302 -2461
rect 265002 -2462 265302 -2461
rect 283002 -2462 283302 -2461
rect 294960 -2462 295260 -2461
rect -3298 -2473 295260 -2462
rect -3298 -2591 -3207 -2473
rect -3089 -2591 13093 -2473
rect 13211 -2591 31093 -2473
rect 31211 -2591 49093 -2473
rect 49211 -2591 67093 -2473
rect 67211 -2591 85093 -2473
rect 85211 -2591 103093 -2473
rect 103211 -2591 121093 -2473
rect 121211 -2591 139093 -2473
rect 139211 -2591 157093 -2473
rect 157211 -2591 175093 -2473
rect 175211 -2591 193093 -2473
rect 193211 -2591 211093 -2473
rect 211211 -2591 229093 -2473
rect 229211 -2591 247093 -2473
rect 247211 -2591 265093 -2473
rect 265211 -2591 283093 -2473
rect 283211 -2591 295051 -2473
rect 295169 -2591 295260 -2473
rect -3298 -2633 295260 -2591
rect -3298 -2751 -3207 -2633
rect -3089 -2751 13093 -2633
rect 13211 -2751 31093 -2633
rect 31211 -2751 49093 -2633
rect 49211 -2751 67093 -2633
rect 67211 -2751 85093 -2633
rect 85211 -2751 103093 -2633
rect 103211 -2751 121093 -2633
rect 121211 -2751 139093 -2633
rect 139211 -2751 157093 -2633
rect 157211 -2751 175093 -2633
rect 175211 -2751 193093 -2633
rect 193211 -2751 211093 -2633
rect 211211 -2751 229093 -2633
rect 229211 -2751 247093 -2633
rect 247211 -2751 265093 -2633
rect 265211 -2751 283093 -2633
rect 283211 -2751 295051 -2633
rect 295169 -2751 295260 -2633
rect -3298 -2762 295260 -2751
rect -3298 -2763 -2998 -2762
rect 13002 -2763 13302 -2762
rect 31002 -2763 31302 -2762
rect 49002 -2763 49302 -2762
rect 67002 -2763 67302 -2762
rect 85002 -2763 85302 -2762
rect 103002 -2763 103302 -2762
rect 121002 -2763 121302 -2762
rect 139002 -2763 139302 -2762
rect 157002 -2763 157302 -2762
rect 175002 -2763 175302 -2762
rect 193002 -2763 193302 -2762
rect 211002 -2763 211302 -2762
rect 229002 -2763 229302 -2762
rect 247002 -2763 247302 -2762
rect 265002 -2763 265302 -2762
rect 283002 -2763 283302 -2762
rect 294960 -2763 295260 -2762
rect -3758 -2922 -3458 -2921
rect 5802 -2922 6102 -2921
rect 23802 -2922 24102 -2921
rect 41802 -2922 42102 -2921
rect 59802 -2922 60102 -2921
rect 77802 -2922 78102 -2921
rect 95802 -2922 96102 -2921
rect 113802 -2922 114102 -2921
rect 131802 -2922 132102 -2921
rect 149802 -2922 150102 -2921
rect 167802 -2922 168102 -2921
rect 185802 -2922 186102 -2921
rect 203802 -2922 204102 -2921
rect 221802 -2922 222102 -2921
rect 239802 -2922 240102 -2921
rect 257802 -2922 258102 -2921
rect 275802 -2922 276102 -2921
rect 295420 -2922 295720 -2921
rect -3758 -2933 295720 -2922
rect -3758 -3051 -3667 -2933
rect -3549 -3051 5893 -2933
rect 6011 -3051 23893 -2933
rect 24011 -3051 41893 -2933
rect 42011 -3051 59893 -2933
rect 60011 -3051 77893 -2933
rect 78011 -3051 95893 -2933
rect 96011 -3051 113893 -2933
rect 114011 -3051 131893 -2933
rect 132011 -3051 149893 -2933
rect 150011 -3051 167893 -2933
rect 168011 -3051 185893 -2933
rect 186011 -3051 203893 -2933
rect 204011 -3051 221893 -2933
rect 222011 -3051 239893 -2933
rect 240011 -3051 257893 -2933
rect 258011 -3051 275893 -2933
rect 276011 -3051 295511 -2933
rect 295629 -3051 295720 -2933
rect -3758 -3093 295720 -3051
rect -3758 -3211 -3667 -3093
rect -3549 -3211 5893 -3093
rect 6011 -3211 23893 -3093
rect 24011 -3211 41893 -3093
rect 42011 -3211 59893 -3093
rect 60011 -3211 77893 -3093
rect 78011 -3211 95893 -3093
rect 96011 -3211 113893 -3093
rect 114011 -3211 131893 -3093
rect 132011 -3211 149893 -3093
rect 150011 -3211 167893 -3093
rect 168011 -3211 185893 -3093
rect 186011 -3211 203893 -3093
rect 204011 -3211 221893 -3093
rect 222011 -3211 239893 -3093
rect 240011 -3211 257893 -3093
rect 258011 -3211 275893 -3093
rect 276011 -3211 295511 -3093
rect 295629 -3211 295720 -3093
rect -3758 -3222 295720 -3211
rect -3758 -3223 -3458 -3222
rect 5802 -3223 6102 -3222
rect 23802 -3223 24102 -3222
rect 41802 -3223 42102 -3222
rect 59802 -3223 60102 -3222
rect 77802 -3223 78102 -3222
rect 95802 -3223 96102 -3222
rect 113802 -3223 114102 -3222
rect 131802 -3223 132102 -3222
rect 149802 -3223 150102 -3222
rect 167802 -3223 168102 -3222
rect 185802 -3223 186102 -3222
rect 203802 -3223 204102 -3222
rect 221802 -3223 222102 -3222
rect 239802 -3223 240102 -3222
rect 257802 -3223 258102 -3222
rect 275802 -3223 276102 -3222
rect 295420 -3223 295720 -3222
rect -4218 -3382 -3918 -3381
rect 14802 -3382 15102 -3381
rect 32802 -3382 33102 -3381
rect 50802 -3382 51102 -3381
rect 68802 -3382 69102 -3381
rect 86802 -3382 87102 -3381
rect 104802 -3382 105102 -3381
rect 122802 -3382 123102 -3381
rect 140802 -3382 141102 -3381
rect 158802 -3382 159102 -3381
rect 176802 -3382 177102 -3381
rect 194802 -3382 195102 -3381
rect 212802 -3382 213102 -3381
rect 230802 -3382 231102 -3381
rect 248802 -3382 249102 -3381
rect 266802 -3382 267102 -3381
rect 284802 -3382 285102 -3381
rect 295880 -3382 296180 -3381
rect -4218 -3393 296180 -3382
rect -4218 -3511 -4127 -3393
rect -4009 -3511 14893 -3393
rect 15011 -3511 32893 -3393
rect 33011 -3511 50893 -3393
rect 51011 -3511 68893 -3393
rect 69011 -3511 86893 -3393
rect 87011 -3511 104893 -3393
rect 105011 -3511 122893 -3393
rect 123011 -3511 140893 -3393
rect 141011 -3511 158893 -3393
rect 159011 -3511 176893 -3393
rect 177011 -3511 194893 -3393
rect 195011 -3511 212893 -3393
rect 213011 -3511 230893 -3393
rect 231011 -3511 248893 -3393
rect 249011 -3511 266893 -3393
rect 267011 -3511 284893 -3393
rect 285011 -3511 295971 -3393
rect 296089 -3511 296180 -3393
rect -4218 -3553 296180 -3511
rect -4218 -3671 -4127 -3553
rect -4009 -3671 14893 -3553
rect 15011 -3671 32893 -3553
rect 33011 -3671 50893 -3553
rect 51011 -3671 68893 -3553
rect 69011 -3671 86893 -3553
rect 87011 -3671 104893 -3553
rect 105011 -3671 122893 -3553
rect 123011 -3671 140893 -3553
rect 141011 -3671 158893 -3553
rect 159011 -3671 176893 -3553
rect 177011 -3671 194893 -3553
rect 195011 -3671 212893 -3553
rect 213011 -3671 230893 -3553
rect 231011 -3671 248893 -3553
rect 249011 -3671 266893 -3553
rect 267011 -3671 284893 -3553
rect 285011 -3671 295971 -3553
rect 296089 -3671 296180 -3553
rect -4218 -3682 296180 -3671
rect -4218 -3683 -3918 -3682
rect 14802 -3683 15102 -3682
rect 32802 -3683 33102 -3682
rect 50802 -3683 51102 -3682
rect 68802 -3683 69102 -3682
rect 86802 -3683 87102 -3682
rect 104802 -3683 105102 -3682
rect 122802 -3683 123102 -3682
rect 140802 -3683 141102 -3682
rect 158802 -3683 159102 -3682
rect 176802 -3683 177102 -3682
rect 194802 -3683 195102 -3682
rect 212802 -3683 213102 -3682
rect 230802 -3683 231102 -3682
rect 248802 -3683 249102 -3682
rect 266802 -3683 267102 -3682
rect 284802 -3683 285102 -3682
rect 295880 -3683 296180 -3682
>>>>>>> upstream/master
<< labels >>
rlabel metal3 s 291760 2898 292480 3018 4 analog_io[0]
port 1 nsew
rlabel metal3 s 291760 237498 292480 237618 4 analog_io[10]
port 2 nsew
rlabel metal3 s 291760 260958 292480 261078 4 analog_io[11]
port 3 nsew
rlabel metal3 s 291760 284418 292480 284538 4 analog_io[12]
port 4 nsew
rlabel metal3 s 291760 307878 292480 307998 4 analog_io[13]
port 5 nsew
rlabel metal3 s 291760 331338 292480 331458 4 analog_io[14]
port 6 nsew
rlabel metal2 s 287909 351760 287965 352480 4 analog_io[15]
port 7 nsew
rlabel metal2 s 255479 351760 255535 352480 4 analog_io[16]
port 8 nsew
rlabel metal2 s 223049 351760 223105 352480 4 analog_io[17]
port 9 nsew
rlabel metal2 s 190573 351760 190629 352480 4 analog_io[18]
port 10 nsew
rlabel metal2 s 158143 351760 158199 352480 4 analog_io[19]
port 11 nsew
rlabel metal3 s 291760 26358 292480 26478 4 analog_io[1]
port 12 nsew
rlabel metal2 s 125713 351760 125769 352480 4 analog_io[20]
port 13 nsew
rlabel metal2 s 93237 351760 93293 352480 4 analog_io[21]
port 14 nsew
rlabel metal2 s 60807 351760 60863 352480 4 analog_io[22]
port 15 nsew
rlabel metal2 s 28377 351760 28433 352480 4 analog_io[23]
port 16 nsew
rlabel metal3 s -480 348270 240 348390 4 analog_io[24]
port 17 nsew
rlabel metal3 s -480 319506 240 319626 4 analog_io[25]
port 18 nsew
rlabel metal3 s -480 290810 240 290930 4 analog_io[26]
port 19 nsew
rlabel metal3 s -480 262046 240 262166 4 analog_io[27]
port 20 nsew
rlabel metal3 s -480 233350 240 233470 4 analog_io[28]
port 21 nsew
rlabel metal3 s -480 204586 240 204706 4 analog_io[29]
port 22 nsew
rlabel metal3 s 291760 49818 292480 49938 4 analog_io[2]
port 23 nsew
rlabel metal3 s -480 175890 240 176010 4 analog_io[30]
port 24 nsew
rlabel metal3 s 291760 73278 292480 73398 4 analog_io[3]
port 25 nsew
rlabel metal3 s 291760 96738 292480 96858 4 analog_io[4]
port 26 nsew
rlabel metal3 s 291760 120198 292480 120318 4 analog_io[5]
port 27 nsew
rlabel metal3 s 291760 143658 292480 143778 4 analog_io[6]
port 28 nsew
rlabel metal3 s 291760 167118 292480 167238 4 analog_io[7]
port 29 nsew
rlabel metal3 s 291760 190578 292480 190698 4 analog_io[8]
port 30 nsew
rlabel metal3 s 291760 214038 292480 214158 4 analog_io[9]
port 31 nsew
rlabel metal3 s 291760 8746 292480 8866 4 io_in[0]
port 32 nsew
rlabel metal3 s 291760 243346 292480 243466 4 io_in[10]
port 33 nsew
rlabel metal3 s 291760 266874 292480 266994 4 io_in[11]
port 34 nsew
rlabel metal3 s 291760 290334 292480 290454 4 io_in[12]
port 35 nsew
rlabel metal3 s 291760 313794 292480 313914 4 io_in[13]
port 36 nsew
rlabel metal3 s 291760 337254 292480 337374 4 io_in[14]
port 37 nsew
rlabel metal2 s 279813 351760 279869 352480 4 io_in[15]
port 38 nsew
rlabel metal2 s 247383 351760 247439 352480 4 io_in[16]
port 39 nsew
rlabel metal2 s 214907 351760 214963 352480 4 io_in[17]
port 40 nsew
rlabel metal2 s 182477 351760 182533 352480 4 io_in[18]
port 41 nsew
rlabel metal2 s 150047 351760 150103 352480 4 io_in[19]
port 42 nsew
rlabel metal3 s 291760 32206 292480 32326 4 io_in[1]
port 43 nsew
rlabel metal2 s 117571 351760 117627 352480 4 io_in[20]
port 44 nsew
rlabel metal2 s 85141 351760 85197 352480 4 io_in[21]
port 45 nsew
rlabel metal2 s 52711 351760 52767 352480 4 io_in[22]
port 46 nsew
rlabel metal2 s 20235 351760 20291 352480 4 io_in[23]
port 47 nsew
rlabel metal3 s -480 341062 240 341182 4 io_in[24]
port 48 nsew
rlabel metal3 s -480 312366 240 312486 4 io_in[25]
port 49 nsew
rlabel metal3 s -480 283602 240 283722 4 io_in[26]
port 50 nsew
rlabel metal3 s -480 254906 240 255026 4 io_in[27]
port 51 nsew
rlabel metal3 s -480 226142 240 226262 4 io_in[28]
port 52 nsew
rlabel metal3 s -480 197446 240 197566 4 io_in[29]
port 53 nsew
rlabel metal3 s 291760 55666 292480 55786 4 io_in[2]
port 54 nsew
rlabel metal3 s -480 168682 240 168802 4 io_in[30]
port 55 nsew
rlabel metal3 s -480 147126 240 147246 4 io_in[31]
port 56 nsew
rlabel metal3 s -480 125570 240 125690 4 io_in[32]
port 57 nsew
rlabel metal3 s -480 104014 240 104134 4 io_in[33]
port 58 nsew
rlabel metal3 s -480 82458 240 82578 4 io_in[34]
port 59 nsew
rlabel metal3 s -480 60970 240 61090 4 io_in[35]
port 60 nsew
rlabel metal3 s -480 39414 240 39534 4 io_in[36]
port 61 nsew
rlabel metal3 s -480 17858 240 17978 4 io_in[37]
port 62 nsew
rlabel metal3 s 291760 79126 292480 79246 4 io_in[3]
port 63 nsew
rlabel metal3 s 291760 102586 292480 102706 4 io_in[4]
port 64 nsew
rlabel metal3 s 291760 126046 292480 126166 4 io_in[5]
port 65 nsew
rlabel metal3 s 291760 149506 292480 149626 4 io_in[6]
port 66 nsew
rlabel metal3 s 291760 172966 292480 173086 4 io_in[7]
port 67 nsew
rlabel metal3 s 291760 196426 292480 196546 4 io_in[8]
port 68 nsew
rlabel metal3 s 291760 219886 292480 220006 4 io_in[9]
port 69 nsew
rlabel metal3 s 291760 20442 292480 20562 4 io_oeb[0]
port 70 nsew
rlabel metal3 s 291760 255110 292480 255230 4 io_oeb[10]
port 71 nsew
rlabel metal3 s 291760 278570 292480 278690 4 io_oeb[11]
port 72 nsew
rlabel metal3 s 291760 302030 292480 302150 4 io_oeb[12]
port 73 nsew
rlabel metal3 s 291760 325490 292480 325610 4 io_oeb[13]
port 74 nsew
rlabel metal3 s 291760 348950 292480 349070 4 io_oeb[14]
port 75 nsew
rlabel metal2 s 263575 351760 263631 352480 4 io_oeb[15]
port 76 nsew
rlabel metal2 s 231145 351760 231201 352480 4 io_oeb[16]
port 77 nsew
rlabel metal2 s 198715 351760 198771 352480 4 io_oeb[17]
port 78 nsew
rlabel metal2 s 166239 351760 166295 352480 4 io_oeb[18]
port 79 nsew
rlabel metal2 s 133809 351760 133865 352480 4 io_oeb[19]
port 80 nsew
rlabel metal3 s 291760 43902 292480 44022 4 io_oeb[1]
port 81 nsew
rlabel metal2 s 101379 351760 101435 352480 4 io_oeb[20]
port 82 nsew
rlabel metal2 s 68903 351760 68959 352480 4 io_oeb[21]
port 83 nsew
rlabel metal2 s 36473 351760 36529 352480 4 io_oeb[22]
port 84 nsew
rlabel metal2 s 4043 351760 4099 352480 4 io_oeb[23]
port 85 nsew
rlabel metal3 s -480 326714 240 326834 4 io_oeb[24]
port 86 nsew
rlabel metal3 s -480 297950 240 298070 4 io_oeb[25]
port 87 nsew
rlabel metal3 s -480 269254 240 269374 4 io_oeb[26]
port 88 nsew
rlabel metal3 s -480 240490 240 240610 4 io_oeb[27]
port 89 nsew
rlabel metal3 s -480 211794 240 211914 4 io_oeb[28]
port 90 nsew
rlabel metal3 s -480 183030 240 183150 4 io_oeb[29]
port 91 nsew
rlabel metal3 s 291760 67362 292480 67482 4 io_oeb[2]
port 92 nsew
rlabel metal3 s -480 154334 240 154454 4 io_oeb[30]
port 93 nsew
rlabel metal3 s -480 132778 240 132898 4 io_oeb[31]
port 94 nsew
rlabel metal3 s -480 111222 240 111342 4 io_oeb[32]
port 95 nsew
rlabel metal3 s -480 89666 240 89786 4 io_oeb[33]
port 96 nsew
rlabel metal3 s -480 68110 240 68230 4 io_oeb[34]
port 97 nsew
rlabel metal3 s -480 46554 240 46674 4 io_oeb[35]
port 98 nsew
rlabel metal3 s -480 24998 240 25118 4 io_oeb[36]
port 99 nsew
rlabel metal3 s -480 3510 240 3630 4 io_oeb[37]
port 100 nsew
rlabel metal3 s 291760 90890 292480 91010 4 io_oeb[3]
port 101 nsew
rlabel metal3 s 291760 114350 292480 114470 4 io_oeb[4]
port 102 nsew
rlabel metal3 s 291760 137810 292480 137930 4 io_oeb[5]
port 103 nsew
rlabel metal3 s 291760 161270 292480 161390 4 io_oeb[6]
port 104 nsew
rlabel metal3 s 291760 184730 292480 184850 4 io_oeb[7]
port 105 nsew
rlabel metal3 s 291760 208190 292480 208310 4 io_oeb[8]
port 106 nsew
rlabel metal3 s 291760 231650 292480 231770 4 io_oeb[9]
port 107 nsew
rlabel metal3 s 291760 14594 292480 14714 4 io_out[0]
port 108 nsew
rlabel metal3 s 291760 249262 292480 249382 4 io_out[10]
port 109 nsew
rlabel metal3 s 291760 272722 292480 272842 4 io_out[11]
port 110 nsew
rlabel metal3 s 291760 296182 292480 296302 4 io_out[12]
port 111 nsew
rlabel metal3 s 291760 319642 292480 319762 4 io_out[13]
port 112 nsew
rlabel metal3 s 291760 343102 292480 343222 4 io_out[14]
port 113 nsew
rlabel metal2 s 271717 351760 271773 352480 4 io_out[15]
port 114 nsew
rlabel metal2 s 239241 351760 239297 352480 4 io_out[16]
port 115 nsew
rlabel metal2 s 206811 351760 206867 352480 4 io_out[17]
port 116 nsew
rlabel metal2 s 174381 351760 174437 352480 4 io_out[18]
port 117 nsew
rlabel metal2 s 141905 351760 141961 352480 4 io_out[19]
port 118 nsew
rlabel metal3 s 291760 38054 292480 38174 4 io_out[1]
port 119 nsew
rlabel metal2 s 109475 351760 109531 352480 4 io_out[20]
port 120 nsew
rlabel metal2 s 77045 351760 77101 352480 4 io_out[21]
port 121 nsew
rlabel metal2 s 44569 351760 44625 352480 4 io_out[22]
port 122 nsew
rlabel metal2 s 12139 351760 12195 352480 4 io_out[23]
port 123 nsew
rlabel metal3 s -480 333922 240 334042 4 io_out[24]
port 124 nsew
rlabel metal3 s -480 305158 240 305278 4 io_out[25]
port 125 nsew
rlabel metal3 s -480 276462 240 276582 4 io_out[26]
port 126 nsew
rlabel metal3 s -480 247698 240 247818 4 io_out[27]
port 127 nsew
rlabel metal3 s -480 218934 240 219054 4 io_out[28]
port 128 nsew
rlabel metal3 s -480 190238 240 190358 4 io_out[29]
port 129 nsew
rlabel metal3 s 291760 61514 292480 61634 4 io_out[2]
port 130 nsew
rlabel metal3 s -480 161474 240 161594 4 io_out[30]
port 131 nsew
rlabel metal3 s -480 139986 240 140106 4 io_out[31]
port 132 nsew
rlabel metal3 s -480 118430 240 118550 4 io_out[32]
port 133 nsew
rlabel metal3 s -480 96874 240 96994 4 io_out[33]
port 134 nsew
rlabel metal3 s -480 75318 240 75438 4 io_out[34]
port 135 nsew
rlabel metal3 s -480 53762 240 53882 4 io_out[35]
port 136 nsew
rlabel metal3 s -480 32206 240 32326 4 io_out[36]
port 137 nsew
rlabel metal3 s -480 10650 240 10770 4 io_out[37]
port 138 nsew
rlabel metal3 s 291760 84974 292480 85094 4 io_out[3]
port 139 nsew
rlabel metal3 s 291760 108434 292480 108554 4 io_out[4]
port 140 nsew
rlabel metal3 s 291760 131894 292480 132014 4 io_out[5]
port 141 nsew
rlabel metal3 s 291760 155354 292480 155474 4 io_out[6]
port 142 nsew
rlabel metal3 s 291760 178882 292480 179002 4 io_out[7]
port 143 nsew
rlabel metal3 s 291760 202342 292480 202462 4 io_out[8]
port 144 nsew
rlabel metal3 s 291760 225802 292480 225922 4 io_out[9]
port 145 nsew
rlabel metal2 s 63291 -480 63347 240 4 la_data_in[0]
port 146 nsew
rlabel metal2 s 241725 -480 241781 240 4 la_data_in[100]
port 147 nsew
rlabel metal2 s 243473 -480 243529 240 4 la_data_in[101]
port 148 nsew
rlabel metal2 s 245267 -480 245323 240 4 la_data_in[102]
port 149 nsew
rlabel metal2 s 247061 -480 247117 240 4 la_data_in[103]
port 150 nsew
rlabel metal2 s 248855 -480 248911 240 4 la_data_in[104]
port 151 nsew
rlabel metal2 s 250603 -480 250659 240 4 la_data_in[105]
port 152 nsew
rlabel metal2 s 252397 -480 252453 240 4 la_data_in[106]
port 153 nsew
rlabel metal2 s 254191 -480 254247 240 4 la_data_in[107]
port 154 nsew
rlabel metal2 s 255985 -480 256041 240 4 la_data_in[108]
port 155 nsew
rlabel metal2 s 257779 -480 257835 240 4 la_data_in[109]
port 156 nsew
rlabel metal2 s 81139 -480 81195 240 4 la_data_in[10]
port 157 nsew
rlabel metal2 s 259527 -480 259583 240 4 la_data_in[110]
port 158 nsew
rlabel metal2 s 261321 -480 261377 240 4 la_data_in[111]
port 159 nsew
rlabel metal2 s 263115 -480 263171 240 4 la_data_in[112]
port 160 nsew
rlabel metal2 s 264909 -480 264965 240 4 la_data_in[113]
port 161 nsew
rlabel metal2 s 266703 -480 266759 240 4 la_data_in[114]
port 162 nsew
rlabel metal2 s 268451 -480 268507 240 4 la_data_in[115]
port 163 nsew
rlabel metal2 s 270245 -480 270301 240 4 la_data_in[116]
port 164 nsew
rlabel metal2 s 272039 -480 272095 240 4 la_data_in[117]
port 165 nsew
rlabel metal2 s 273833 -480 273889 240 4 la_data_in[118]
port 166 nsew
rlabel metal2 s 275581 -480 275637 240 4 la_data_in[119]
port 167 nsew
rlabel metal2 s 82933 -480 82989 240 4 la_data_in[11]
port 168 nsew
rlabel metal2 s 277375 -480 277431 240 4 la_data_in[120]
port 169 nsew
rlabel metal2 s 279169 -480 279225 240 4 la_data_in[121]
port 170 nsew
rlabel metal2 s 280963 -480 281019 240 4 la_data_in[122]
port 171 nsew
rlabel metal2 s 282757 -480 282813 240 4 la_data_in[123]
port 172 nsew
rlabel metal2 s 284505 -480 284561 240 4 la_data_in[124]
port 173 nsew
rlabel metal2 s 286299 -480 286355 240 4 la_data_in[125]
port 174 nsew
rlabel metal2 s 288093 -480 288149 240 4 la_data_in[126]
port 175 nsew
rlabel metal2 s 289887 -480 289943 240 4 la_data_in[127]
port 176 nsew
rlabel metal2 s 84681 -480 84737 240 4 la_data_in[12]
port 177 nsew
rlabel metal2 s 86475 -480 86531 240 4 la_data_in[13]
port 178 nsew
rlabel metal2 s 88269 -480 88325 240 4 la_data_in[14]
port 179 nsew
rlabel metal2 s 90063 -480 90119 240 4 la_data_in[15]
port 180 nsew
rlabel metal2 s 91857 -480 91913 240 4 la_data_in[16]
port 181 nsew
rlabel metal2 s 93605 -480 93661 240 4 la_data_in[17]
port 182 nsew
rlabel metal2 s 95399 -480 95455 240 4 la_data_in[18]
port 183 nsew
rlabel metal2 s 97193 -480 97249 240 4 la_data_in[19]
port 184 nsew
rlabel metal2 s 65085 -480 65141 240 4 la_data_in[1]
port 185 nsew
rlabel metal2 s 98987 -480 99043 240 4 la_data_in[20]
port 186 nsew
rlabel metal2 s 100735 -480 100791 240 4 la_data_in[21]
port 187 nsew
rlabel metal2 s 102529 -480 102585 240 4 la_data_in[22]
port 188 nsew
rlabel metal2 s 104323 -480 104379 240 4 la_data_in[23]
port 189 nsew
rlabel metal2 s 106117 -480 106173 240 4 la_data_in[24]
port 190 nsew
rlabel metal2 s 107911 -480 107967 240 4 la_data_in[25]
port 191 nsew
rlabel metal2 s 109659 -480 109715 240 4 la_data_in[26]
port 192 nsew
rlabel metal2 s 111453 -480 111509 240 4 la_data_in[27]
port 193 nsew
rlabel metal2 s 113247 -480 113303 240 4 la_data_in[28]
port 194 nsew
rlabel metal2 s 115041 -480 115097 240 4 la_data_in[29]
port 195 nsew
rlabel metal2 s 66879 -480 66935 240 4 la_data_in[2]
port 196 nsew
rlabel metal2 s 116835 -480 116891 240 4 la_data_in[30]
port 197 nsew
rlabel metal2 s 118583 -480 118639 240 4 la_data_in[31]
port 198 nsew
rlabel metal2 s 120377 -480 120433 240 4 la_data_in[32]
port 199 nsew
rlabel metal2 s 122171 -480 122227 240 4 la_data_in[33]
port 200 nsew
rlabel metal2 s 123965 -480 124021 240 4 la_data_in[34]
port 201 nsew
rlabel metal2 s 125713 -480 125769 240 4 la_data_in[35]
port 202 nsew
rlabel metal2 s 127507 -480 127563 240 4 la_data_in[36]
port 203 nsew
rlabel metal2 s 129301 -480 129357 240 4 la_data_in[37]
port 204 nsew
rlabel metal2 s 131095 -480 131151 240 4 la_data_in[38]
port 205 nsew
rlabel metal2 s 132889 -480 132945 240 4 la_data_in[39]
port 206 nsew
rlabel metal2 s 68627 -480 68683 240 4 la_data_in[3]
port 207 nsew
rlabel metal2 s 134637 -480 134693 240 4 la_data_in[40]
port 208 nsew
rlabel metal2 s 136431 -480 136487 240 4 la_data_in[41]
port 209 nsew
rlabel metal2 s 138225 -480 138281 240 4 la_data_in[42]
port 210 nsew
rlabel metal2 s 140019 -480 140075 240 4 la_data_in[43]
port 211 nsew
rlabel metal2 s 141813 -480 141869 240 4 la_data_in[44]
port 212 nsew
rlabel metal2 s 143561 -480 143617 240 4 la_data_in[45]
port 213 nsew
rlabel metal2 s 145355 -480 145411 240 4 la_data_in[46]
port 214 nsew
rlabel metal2 s 147149 -480 147205 240 4 la_data_in[47]
port 215 nsew
rlabel metal2 s 148943 -480 148999 240 4 la_data_in[48]
port 216 nsew
rlabel metal2 s 150691 -480 150747 240 4 la_data_in[49]
port 217 nsew
rlabel metal2 s 70421 -480 70477 240 4 la_data_in[4]
port 218 nsew
rlabel metal2 s 152485 -480 152541 240 4 la_data_in[50]
port 219 nsew
rlabel metal2 s 154279 -480 154335 240 4 la_data_in[51]
port 220 nsew
rlabel metal2 s 156073 -480 156129 240 4 la_data_in[52]
port 221 nsew
rlabel metal2 s 157867 -480 157923 240 4 la_data_in[53]
port 222 nsew
rlabel metal2 s 159615 -480 159671 240 4 la_data_in[54]
port 223 nsew
rlabel metal2 s 161409 -480 161465 240 4 la_data_in[55]
port 224 nsew
rlabel metal2 s 163203 -480 163259 240 4 la_data_in[56]
port 225 nsew
rlabel metal2 s 164997 -480 165053 240 4 la_data_in[57]
port 226 nsew
rlabel metal2 s 166791 -480 166847 240 4 la_data_in[58]
port 227 nsew
rlabel metal2 s 168539 -480 168595 240 4 la_data_in[59]
port 228 nsew
rlabel metal2 s 72215 -480 72271 240 4 la_data_in[5]
port 229 nsew
rlabel metal2 s 170333 -480 170389 240 4 la_data_in[60]
port 230 nsew
rlabel metal2 s 172127 -480 172183 240 4 la_data_in[61]
port 231 nsew
rlabel metal2 s 173921 -480 173977 240 4 la_data_in[62]
port 232 nsew
rlabel metal2 s 175669 -480 175725 240 4 la_data_in[63]
port 233 nsew
rlabel metal2 s 177463 -480 177519 240 4 la_data_in[64]
port 234 nsew
rlabel metal2 s 179257 -480 179313 240 4 la_data_in[65]
port 235 nsew
rlabel metal2 s 181051 -480 181107 240 4 la_data_in[66]
port 236 nsew
rlabel metal2 s 182845 -480 182901 240 4 la_data_in[67]
port 237 nsew
rlabel metal2 s 184593 -480 184649 240 4 la_data_in[68]
port 238 nsew
rlabel metal2 s 186387 -480 186443 240 4 la_data_in[69]
port 239 nsew
rlabel metal2 s 74009 -480 74065 240 4 la_data_in[6]
port 240 nsew
rlabel metal2 s 188181 -480 188237 240 4 la_data_in[70]
port 241 nsew
rlabel metal2 s 189975 -480 190031 240 4 la_data_in[71]
port 242 nsew
rlabel metal2 s 191769 -480 191825 240 4 la_data_in[72]
port 243 nsew
rlabel metal2 s 193517 -480 193573 240 4 la_data_in[73]
port 244 nsew
rlabel metal2 s 195311 -480 195367 240 4 la_data_in[74]
port 245 nsew
rlabel metal2 s 197105 -480 197161 240 4 la_data_in[75]
port 246 nsew
rlabel metal2 s 198899 -480 198955 240 4 la_data_in[76]
port 247 nsew
rlabel metal2 s 200647 -480 200703 240 4 la_data_in[77]
port 248 nsew
rlabel metal2 s 202441 -480 202497 240 4 la_data_in[78]
port 249 nsew
rlabel metal2 s 204235 -480 204291 240 4 la_data_in[79]
port 250 nsew
rlabel metal2 s 75757 -480 75813 240 4 la_data_in[7]
port 251 nsew
rlabel metal2 s 206029 -480 206085 240 4 la_data_in[80]
port 252 nsew
rlabel metal2 s 207823 -480 207879 240 4 la_data_in[81]
port 253 nsew
rlabel metal2 s 209571 -480 209627 240 4 la_data_in[82]
port 254 nsew
rlabel metal2 s 211365 -480 211421 240 4 la_data_in[83]
port 255 nsew
rlabel metal2 s 213159 -480 213215 240 4 la_data_in[84]
port 256 nsew
rlabel metal2 s 214953 -480 215009 240 4 la_data_in[85]
port 257 nsew
rlabel metal2 s 216747 -480 216803 240 4 la_data_in[86]
port 258 nsew
rlabel metal2 s 218495 -480 218551 240 4 la_data_in[87]
port 259 nsew
rlabel metal2 s 220289 -480 220345 240 4 la_data_in[88]
port 260 nsew
rlabel metal2 s 222083 -480 222139 240 4 la_data_in[89]
port 261 nsew
rlabel metal2 s 77551 -480 77607 240 4 la_data_in[8]
port 262 nsew
rlabel metal2 s 223877 -480 223933 240 4 la_data_in[90]
port 263 nsew
rlabel metal2 s 225625 -480 225681 240 4 la_data_in[91]
port 264 nsew
rlabel metal2 s 227419 -480 227475 240 4 la_data_in[92]
port 265 nsew
rlabel metal2 s 229213 -480 229269 240 4 la_data_in[93]
port 266 nsew
rlabel metal2 s 231007 -480 231063 240 4 la_data_in[94]
port 267 nsew
rlabel metal2 s 232801 -480 232857 240 4 la_data_in[95]
port 268 nsew
rlabel metal2 s 234549 -480 234605 240 4 la_data_in[96]
port 269 nsew
rlabel metal2 s 236343 -480 236399 240 4 la_data_in[97]
port 270 nsew
rlabel metal2 s 238137 -480 238193 240 4 la_data_in[98]
port 271 nsew
rlabel metal2 s 239931 -480 239987 240 4 la_data_in[99]
port 272 nsew
rlabel metal2 s 79345 -480 79401 240 4 la_data_in[9]
port 273 nsew
rlabel metal2 s 63889 -480 63945 240 4 la_data_out[0]
port 274 nsew
rlabel metal2 s 242277 -480 242333 240 4 la_data_out[100]
port 275 nsew
rlabel metal2 s 244071 -480 244127 240 4 la_data_out[101]
port 276 nsew
rlabel metal2 s 245865 -480 245921 240 4 la_data_out[102]
port 277 nsew
rlabel metal2 s 247659 -480 247715 240 4 la_data_out[103]
port 278 nsew
rlabel metal2 s 249453 -480 249509 240 4 la_data_out[104]
port 279 nsew
rlabel metal2 s 251201 -480 251257 240 4 la_data_out[105]
port 280 nsew
rlabel metal2 s 252995 -480 253051 240 4 la_data_out[106]
port 281 nsew
rlabel metal2 s 254789 -480 254845 240 4 la_data_out[107]
port 282 nsew
rlabel metal2 s 256583 -480 256639 240 4 la_data_out[108]
port 283 nsew
rlabel metal2 s 258377 -480 258433 240 4 la_data_out[109]
port 284 nsew
rlabel metal2 s 81737 -480 81793 240 4 la_data_out[10]
port 285 nsew
rlabel metal2 s 260125 -480 260181 240 4 la_data_out[110]
port 286 nsew
rlabel metal2 s 261919 -480 261975 240 4 la_data_out[111]
port 287 nsew
rlabel metal2 s 263713 -480 263769 240 4 la_data_out[112]
port 288 nsew
rlabel metal2 s 265507 -480 265563 240 4 la_data_out[113]
port 289 nsew
rlabel metal2 s 267255 -480 267311 240 4 la_data_out[114]
port 290 nsew
rlabel metal2 s 269049 -480 269105 240 4 la_data_out[115]
port 291 nsew
rlabel metal2 s 270843 -480 270899 240 4 la_data_out[116]
port 292 nsew
rlabel metal2 s 272637 -480 272693 240 4 la_data_out[117]
port 293 nsew
rlabel metal2 s 274431 -480 274487 240 4 la_data_out[118]
port 294 nsew
rlabel metal2 s 276179 -480 276235 240 4 la_data_out[119]
port 295 nsew
rlabel metal2 s 83531 -480 83587 240 4 la_data_out[11]
port 296 nsew
rlabel metal2 s 277973 -480 278029 240 4 la_data_out[120]
port 297 nsew
rlabel metal2 s 279767 -480 279823 240 4 la_data_out[121]
port 298 nsew
rlabel metal2 s 281561 -480 281617 240 4 la_data_out[122]
port 299 nsew
rlabel metal2 s 283355 -480 283411 240 4 la_data_out[123]
port 300 nsew
rlabel metal2 s 285103 -480 285159 240 4 la_data_out[124]
port 301 nsew
rlabel metal2 s 286897 -480 286953 240 4 la_data_out[125]
port 302 nsew
rlabel metal2 s 288691 -480 288747 240 4 la_data_out[126]
port 303 nsew
rlabel metal2 s 290485 -480 290541 240 4 la_data_out[127]
port 304 nsew
rlabel metal2 s 85279 -480 85335 240 4 la_data_out[12]
port 305 nsew
rlabel metal2 s 87073 -480 87129 240 4 la_data_out[13]
port 306 nsew
rlabel metal2 s 88867 -480 88923 240 4 la_data_out[14]
port 307 nsew
rlabel metal2 s 90661 -480 90717 240 4 la_data_out[15]
port 308 nsew
rlabel metal2 s 92409 -480 92465 240 4 la_data_out[16]
port 309 nsew
rlabel metal2 s 94203 -480 94259 240 4 la_data_out[17]
port 310 nsew
rlabel metal2 s 95997 -480 96053 240 4 la_data_out[18]
port 311 nsew
rlabel metal2 s 97791 -480 97847 240 4 la_data_out[19]
port 312 nsew
rlabel metal2 s 65683 -480 65739 240 4 la_data_out[1]
port 313 nsew
rlabel metal2 s 99585 -480 99641 240 4 la_data_out[20]
port 314 nsew
rlabel metal2 s 101333 -480 101389 240 4 la_data_out[21]
port 315 nsew
rlabel metal2 s 103127 -480 103183 240 4 la_data_out[22]
port 316 nsew
rlabel metal2 s 104921 -480 104977 240 4 la_data_out[23]
port 317 nsew
rlabel metal2 s 106715 -480 106771 240 4 la_data_out[24]
port 318 nsew
rlabel metal2 s 108509 -480 108565 240 4 la_data_out[25]
port 319 nsew
rlabel metal2 s 110257 -480 110313 240 4 la_data_out[26]
port 320 nsew
rlabel metal2 s 112051 -480 112107 240 4 la_data_out[27]
port 321 nsew
rlabel metal2 s 113845 -480 113901 240 4 la_data_out[28]
port 322 nsew
rlabel metal2 s 115639 -480 115695 240 4 la_data_out[29]
port 323 nsew
rlabel metal2 s 67431 -480 67487 240 4 la_data_out[2]
port 324 nsew
rlabel metal2 s 117387 -480 117443 240 4 la_data_out[30]
port 325 nsew
rlabel metal2 s 119181 -480 119237 240 4 la_data_out[31]
port 326 nsew
rlabel metal2 s 120975 -480 121031 240 4 la_data_out[32]
port 327 nsew
rlabel metal2 s 122769 -480 122825 240 4 la_data_out[33]
port 328 nsew
rlabel metal2 s 124563 -480 124619 240 4 la_data_out[34]
port 329 nsew
rlabel metal2 s 126311 -480 126367 240 4 la_data_out[35]
port 330 nsew
rlabel metal2 s 128105 -480 128161 240 4 la_data_out[36]
port 331 nsew
rlabel metal2 s 129899 -480 129955 240 4 la_data_out[37]
port 332 nsew
rlabel metal2 s 131693 -480 131749 240 4 la_data_out[38]
port 333 nsew
rlabel metal2 s 133487 -480 133543 240 4 la_data_out[39]
port 334 nsew
rlabel metal2 s 69225 -480 69281 240 4 la_data_out[3]
port 335 nsew
rlabel metal2 s 135235 -480 135291 240 4 la_data_out[40]
port 336 nsew
rlabel metal2 s 137029 -480 137085 240 4 la_data_out[41]
port 337 nsew
rlabel metal2 s 138823 -480 138879 240 4 la_data_out[42]
port 338 nsew
rlabel metal2 s 140617 -480 140673 240 4 la_data_out[43]
port 339 nsew
rlabel metal2 s 142365 -480 142421 240 4 la_data_out[44]
port 340 nsew
rlabel metal2 s 144159 -480 144215 240 4 la_data_out[45]
port 341 nsew
rlabel metal2 s 145953 -480 146009 240 4 la_data_out[46]
port 342 nsew
rlabel metal2 s 147747 -480 147803 240 4 la_data_out[47]
port 343 nsew
rlabel metal2 s 149541 -480 149597 240 4 la_data_out[48]
port 344 nsew
rlabel metal2 s 151289 -480 151345 240 4 la_data_out[49]
port 345 nsew
rlabel metal2 s 71019 -480 71075 240 4 la_data_out[4]
port 346 nsew
rlabel metal2 s 153083 -480 153139 240 4 la_data_out[50]
port 347 nsew
rlabel metal2 s 154877 -480 154933 240 4 la_data_out[51]
port 348 nsew
rlabel metal2 s 156671 -480 156727 240 4 la_data_out[52]
port 349 nsew
rlabel metal2 s 158465 -480 158521 240 4 la_data_out[53]
port 350 nsew
rlabel metal2 s 160213 -480 160269 240 4 la_data_out[54]
port 351 nsew
rlabel metal2 s 162007 -480 162063 240 4 la_data_out[55]
port 352 nsew
rlabel metal2 s 163801 -480 163857 240 4 la_data_out[56]
port 353 nsew
rlabel metal2 s 165595 -480 165651 240 4 la_data_out[57]
port 354 nsew
rlabel metal2 s 167343 -480 167399 240 4 la_data_out[58]
port 355 nsew
rlabel metal2 s 169137 -480 169193 240 4 la_data_out[59]
port 356 nsew
rlabel metal2 s 72813 -480 72869 240 4 la_data_out[5]
port 357 nsew
rlabel metal2 s 170931 -480 170987 240 4 la_data_out[60]
port 358 nsew
rlabel metal2 s 172725 -480 172781 240 4 la_data_out[61]
port 359 nsew
rlabel metal2 s 174519 -480 174575 240 4 la_data_out[62]
port 360 nsew
rlabel metal2 s 176267 -480 176323 240 4 la_data_out[63]
port 361 nsew
rlabel metal2 s 178061 -480 178117 240 4 la_data_out[64]
port 362 nsew
rlabel metal2 s 179855 -480 179911 240 4 la_data_out[65]
port 363 nsew
rlabel metal2 s 181649 -480 181705 240 4 la_data_out[66]
port 364 nsew
rlabel metal2 s 183443 -480 183499 240 4 la_data_out[67]
port 365 nsew
rlabel metal2 s 185191 -480 185247 240 4 la_data_out[68]
port 366 nsew
rlabel metal2 s 186985 -480 187041 240 4 la_data_out[69]
port 367 nsew
rlabel metal2 s 74607 -480 74663 240 4 la_data_out[6]
port 368 nsew
rlabel metal2 s 188779 -480 188835 240 4 la_data_out[70]
port 369 nsew
rlabel metal2 s 190573 -480 190629 240 4 la_data_out[71]
port 370 nsew
rlabel metal2 s 192321 -480 192377 240 4 la_data_out[72]
port 371 nsew
rlabel metal2 s 194115 -480 194171 240 4 la_data_out[73]
port 372 nsew
rlabel metal2 s 195909 -480 195965 240 4 la_data_out[74]
port 373 nsew
rlabel metal2 s 197703 -480 197759 240 4 la_data_out[75]
port 374 nsew
rlabel metal2 s 199497 -480 199553 240 4 la_data_out[76]
port 375 nsew
rlabel metal2 s 201245 -480 201301 240 4 la_data_out[77]
port 376 nsew
rlabel metal2 s 203039 -480 203095 240 4 la_data_out[78]
port 377 nsew
rlabel metal2 s 204833 -480 204889 240 4 la_data_out[79]
port 378 nsew
rlabel metal2 s 76355 -480 76411 240 4 la_data_out[7]
port 379 nsew
rlabel metal2 s 206627 -480 206683 240 4 la_data_out[80]
port 380 nsew
rlabel metal2 s 208421 -480 208477 240 4 la_data_out[81]
port 381 nsew
rlabel metal2 s 210169 -480 210225 240 4 la_data_out[82]
port 382 nsew
rlabel metal2 s 211963 -480 212019 240 4 la_data_out[83]
port 383 nsew
rlabel metal2 s 213757 -480 213813 240 4 la_data_out[84]
port 384 nsew
rlabel metal2 s 215551 -480 215607 240 4 la_data_out[85]
port 385 nsew
rlabel metal2 s 217299 -480 217355 240 4 la_data_out[86]
port 386 nsew
rlabel metal2 s 219093 -480 219149 240 4 la_data_out[87]
port 387 nsew
rlabel metal2 s 220887 -480 220943 240 4 la_data_out[88]
port 388 nsew
rlabel metal2 s 222681 -480 222737 240 4 la_data_out[89]
port 389 nsew
rlabel metal2 s 78149 -480 78205 240 4 la_data_out[8]
port 390 nsew
rlabel metal2 s 224475 -480 224531 240 4 la_data_out[90]
port 391 nsew
rlabel metal2 s 226223 -480 226279 240 4 la_data_out[91]
port 392 nsew
rlabel metal2 s 228017 -480 228073 240 4 la_data_out[92]
port 393 nsew
rlabel metal2 s 229811 -480 229867 240 4 la_data_out[93]
port 394 nsew
rlabel metal2 s 231605 -480 231661 240 4 la_data_out[94]
port 395 nsew
rlabel metal2 s 233399 -480 233455 240 4 la_data_out[95]
port 396 nsew
rlabel metal2 s 235147 -480 235203 240 4 la_data_out[96]
port 397 nsew
rlabel metal2 s 236941 -480 236997 240 4 la_data_out[97]
port 398 nsew
rlabel metal2 s 238735 -480 238791 240 4 la_data_out[98]
port 399 nsew
rlabel metal2 s 240529 -480 240585 240 4 la_data_out[99]
port 400 nsew
rlabel metal2 s 79943 -480 79999 240 4 la_data_out[9]
port 401 nsew
rlabel metal2 s 64487 -480 64543 240 4 la_oen[0]
port 402 nsew
rlabel metal2 s 242875 -480 242931 240 4 la_oen[100]
port 403 nsew
rlabel metal2 s 244669 -480 244725 240 4 la_oen[101]
port 404 nsew
rlabel metal2 s 246463 -480 246519 240 4 la_oen[102]
port 405 nsew
rlabel metal2 s 248257 -480 248313 240 4 la_oen[103]
port 406 nsew
rlabel metal2 s 250051 -480 250107 240 4 la_oen[104]
port 407 nsew
rlabel metal2 s 251799 -480 251855 240 4 la_oen[105]
port 408 nsew
rlabel metal2 s 253593 -480 253649 240 4 la_oen[106]
port 409 nsew
rlabel metal2 s 255387 -480 255443 240 4 la_oen[107]
port 410 nsew
rlabel metal2 s 257181 -480 257237 240 4 la_oen[108]
port 411 nsew
rlabel metal2 s 258929 -480 258985 240 4 la_oen[109]
port 412 nsew
rlabel metal2 s 82335 -480 82391 240 4 la_oen[10]
port 413 nsew
rlabel metal2 s 260723 -480 260779 240 4 la_oen[110]
port 414 nsew
rlabel metal2 s 262517 -480 262573 240 4 la_oen[111]
port 415 nsew
rlabel metal2 s 264311 -480 264367 240 4 la_oen[112]
port 416 nsew
rlabel metal2 s 266105 -480 266161 240 4 la_oen[113]
port 417 nsew
rlabel metal2 s 267853 -480 267909 240 4 la_oen[114]
port 418 nsew
rlabel metal2 s 269647 -480 269703 240 4 la_oen[115]
port 419 nsew
rlabel metal2 s 271441 -480 271497 240 4 la_oen[116]
port 420 nsew
rlabel metal2 s 273235 -480 273291 240 4 la_oen[117]
port 421 nsew
rlabel metal2 s 275029 -480 275085 240 4 la_oen[118]
port 422 nsew
rlabel metal2 s 276777 -480 276833 240 4 la_oen[119]
port 423 nsew
rlabel metal2 s 84083 -480 84139 240 4 la_oen[11]
port 424 nsew
rlabel metal2 s 278571 -480 278627 240 4 la_oen[120]
port 425 nsew
rlabel metal2 s 280365 -480 280421 240 4 la_oen[121]
port 426 nsew
rlabel metal2 s 282159 -480 282215 240 4 la_oen[122]
port 427 nsew
rlabel metal2 s 283907 -480 283963 240 4 la_oen[123]
port 428 nsew
rlabel metal2 s 285701 -480 285757 240 4 la_oen[124]
port 429 nsew
rlabel metal2 s 287495 -480 287551 240 4 la_oen[125]
port 430 nsew
rlabel metal2 s 289289 -480 289345 240 4 la_oen[126]
port 431 nsew
rlabel metal2 s 291083 -480 291139 240 4 la_oen[127]
port 432 nsew
rlabel metal2 s 85877 -480 85933 240 4 la_oen[12]
port 433 nsew
rlabel metal2 s 87671 -480 87727 240 4 la_oen[13]
port 434 nsew
rlabel metal2 s 89465 -480 89521 240 4 la_oen[14]
port 435 nsew
rlabel metal2 s 91259 -480 91315 240 4 la_oen[15]
port 436 nsew
rlabel metal2 s 93007 -480 93063 240 4 la_oen[16]
port 437 nsew
rlabel metal2 s 94801 -480 94857 240 4 la_oen[17]
port 438 nsew
rlabel metal2 s 96595 -480 96651 240 4 la_oen[18]
port 439 nsew
rlabel metal2 s 98389 -480 98445 240 4 la_oen[19]
port 440 nsew
rlabel metal2 s 66281 -480 66337 240 4 la_oen[1]
port 441 nsew
rlabel metal2 s 100183 -480 100239 240 4 la_oen[20]
port 442 nsew
rlabel metal2 s 101931 -480 101987 240 4 la_oen[21]
port 443 nsew
rlabel metal2 s 103725 -480 103781 240 4 la_oen[22]
port 444 nsew
rlabel metal2 s 105519 -480 105575 240 4 la_oen[23]
port 445 nsew
rlabel metal2 s 107313 -480 107369 240 4 la_oen[24]
port 446 nsew
rlabel metal2 s 109061 -480 109117 240 4 la_oen[25]
port 447 nsew
rlabel metal2 s 110855 -480 110911 240 4 la_oen[26]
port 448 nsew
rlabel metal2 s 112649 -480 112705 240 4 la_oen[27]
port 449 nsew
rlabel metal2 s 114443 -480 114499 240 4 la_oen[28]
port 450 nsew
rlabel metal2 s 116237 -480 116293 240 4 la_oen[29]
port 451 nsew
rlabel metal2 s 68029 -480 68085 240 4 la_oen[2]
port 452 nsew
rlabel metal2 s 117985 -480 118041 240 4 la_oen[30]
port 453 nsew
rlabel metal2 s 119779 -480 119835 240 4 la_oen[31]
port 454 nsew
rlabel metal2 s 121573 -480 121629 240 4 la_oen[32]
port 455 nsew
rlabel metal2 s 123367 -480 123423 240 4 la_oen[33]
port 456 nsew
rlabel metal2 s 125161 -480 125217 240 4 la_oen[34]
port 457 nsew
rlabel metal2 s 126909 -480 126965 240 4 la_oen[35]
port 458 nsew
rlabel metal2 s 128703 -480 128759 240 4 la_oen[36]
port 459 nsew
rlabel metal2 s 130497 -480 130553 240 4 la_oen[37]
port 460 nsew
rlabel metal2 s 132291 -480 132347 240 4 la_oen[38]
port 461 nsew
rlabel metal2 s 134039 -480 134095 240 4 la_oen[39]
port 462 nsew
rlabel metal2 s 69823 -480 69879 240 4 la_oen[3]
port 463 nsew
rlabel metal2 s 135833 -480 135889 240 4 la_oen[40]
port 464 nsew
rlabel metal2 s 137627 -480 137683 240 4 la_oen[41]
port 465 nsew
rlabel metal2 s 139421 -480 139477 240 4 la_oen[42]
port 466 nsew
rlabel metal2 s 141215 -480 141271 240 4 la_oen[43]
port 467 nsew
rlabel metal2 s 142963 -480 143019 240 4 la_oen[44]
port 468 nsew
rlabel metal2 s 144757 -480 144813 240 4 la_oen[45]
port 469 nsew
rlabel metal2 s 146551 -480 146607 240 4 la_oen[46]
port 470 nsew
rlabel metal2 s 148345 -480 148401 240 4 la_oen[47]
port 471 nsew
rlabel metal2 s 150139 -480 150195 240 4 la_oen[48]
port 472 nsew
rlabel metal2 s 151887 -480 151943 240 4 la_oen[49]
port 473 nsew
rlabel metal2 s 71617 -480 71673 240 4 la_oen[4]
port 474 nsew
rlabel metal2 s 153681 -480 153737 240 4 la_oen[50]
port 475 nsew
rlabel metal2 s 155475 -480 155531 240 4 la_oen[51]
port 476 nsew
rlabel metal2 s 157269 -480 157325 240 4 la_oen[52]
port 477 nsew
rlabel metal2 s 159017 -480 159073 240 4 la_oen[53]
port 478 nsew
rlabel metal2 s 160811 -480 160867 240 4 la_oen[54]
port 479 nsew
rlabel metal2 s 162605 -480 162661 240 4 la_oen[55]
port 480 nsew
rlabel metal2 s 164399 -480 164455 240 4 la_oen[56]
port 481 nsew
rlabel metal2 s 166193 -480 166249 240 4 la_oen[57]
port 482 nsew
rlabel metal2 s 167941 -480 167997 240 4 la_oen[58]
port 483 nsew
rlabel metal2 s 169735 -480 169791 240 4 la_oen[59]
port 484 nsew
rlabel metal2 s 73411 -480 73467 240 4 la_oen[5]
port 485 nsew
rlabel metal2 s 171529 -480 171585 240 4 la_oen[60]
port 486 nsew
rlabel metal2 s 173323 -480 173379 240 4 la_oen[61]
port 487 nsew
rlabel metal2 s 175117 -480 175173 240 4 la_oen[62]
port 488 nsew
rlabel metal2 s 176865 -480 176921 240 4 la_oen[63]
port 489 nsew
rlabel metal2 s 178659 -480 178715 240 4 la_oen[64]
port 490 nsew
rlabel metal2 s 180453 -480 180509 240 4 la_oen[65]
port 491 nsew
rlabel metal2 s 182247 -480 182303 240 4 la_oen[66]
port 492 nsew
rlabel metal2 s 183995 -480 184051 240 4 la_oen[67]
port 493 nsew
rlabel metal2 s 185789 -480 185845 240 4 la_oen[68]
port 494 nsew
rlabel metal2 s 187583 -480 187639 240 4 la_oen[69]
port 495 nsew
rlabel metal2 s 75205 -480 75261 240 4 la_oen[6]
port 496 nsew
rlabel metal2 s 189377 -480 189433 240 4 la_oen[70]
port 497 nsew
rlabel metal2 s 191171 -480 191227 240 4 la_oen[71]
port 498 nsew
rlabel metal2 s 192919 -480 192975 240 4 la_oen[72]
port 499 nsew
rlabel metal2 s 194713 -480 194769 240 4 la_oen[73]
port 500 nsew
rlabel metal2 s 196507 -480 196563 240 4 la_oen[74]
port 501 nsew
rlabel metal2 s 198301 -480 198357 240 4 la_oen[75]
port 502 nsew
rlabel metal2 s 200095 -480 200151 240 4 la_oen[76]
port 503 nsew
rlabel metal2 s 201843 -480 201899 240 4 la_oen[77]
port 504 nsew
rlabel metal2 s 203637 -480 203693 240 4 la_oen[78]
port 505 nsew
rlabel metal2 s 205431 -480 205487 240 4 la_oen[79]
port 506 nsew
rlabel metal2 s 76953 -480 77009 240 4 la_oen[7]
port 507 nsew
rlabel metal2 s 207225 -480 207281 240 4 la_oen[80]
port 508 nsew
rlabel metal2 s 208973 -480 209029 240 4 la_oen[81]
port 509 nsew
rlabel metal2 s 210767 -480 210823 240 4 la_oen[82]
port 510 nsew
rlabel metal2 s 212561 -480 212617 240 4 la_oen[83]
port 511 nsew
rlabel metal2 s 214355 -480 214411 240 4 la_oen[84]
port 512 nsew
rlabel metal2 s 216149 -480 216205 240 4 la_oen[85]
port 513 nsew
rlabel metal2 s 217897 -480 217953 240 4 la_oen[86]
port 514 nsew
rlabel metal2 s 219691 -480 219747 240 4 la_oen[87]
port 515 nsew
rlabel metal2 s 221485 -480 221541 240 4 la_oen[88]
port 516 nsew
rlabel metal2 s 223279 -480 223335 240 4 la_oen[89]
port 517 nsew
rlabel metal2 s 78747 -480 78803 240 4 la_oen[8]
port 518 nsew
rlabel metal2 s 225073 -480 225129 240 4 la_oen[90]
port 519 nsew
rlabel metal2 s 226821 -480 226877 240 4 la_oen[91]
port 520 nsew
rlabel metal2 s 228615 -480 228671 240 4 la_oen[92]
port 521 nsew
rlabel metal2 s 230409 -480 230465 240 4 la_oen[93]
port 522 nsew
rlabel metal2 s 232203 -480 232259 240 4 la_oen[94]
port 523 nsew
rlabel metal2 s 233951 -480 234007 240 4 la_oen[95]
port 524 nsew
rlabel metal2 s 235745 -480 235801 240 4 la_oen[96]
port 525 nsew
rlabel metal2 s 237539 -480 237595 240 4 la_oen[97]
port 526 nsew
rlabel metal2 s 239333 -480 239389 240 4 la_oen[98]
port 527 nsew
rlabel metal2 s 241127 -480 241183 240 4 la_oen[99]
port 528 nsew
rlabel metal2 s 80541 -480 80597 240 4 la_oen[9]
port 529 nsew
rlabel metal2 s 291681 -480 291737 240 4 user_clock2
port 530 nsew
rlabel metal2 s 271 -480 327 240 4 wb_clk_i
port 531 nsew
rlabel metal2 s 823 -480 879 240 4 wb_rst_i
port 532 nsew
rlabel metal2 s 1421 -480 1477 240 4 wbs_ack_o
port 533 nsew
rlabel metal2 s 3813 -480 3869 240 4 wbs_adr_i[0]
port 534 nsew
rlabel metal2 s 24053 -480 24109 240 4 wbs_adr_i[10]
port 535 nsew
rlabel metal2 s 25801 -480 25857 240 4 wbs_adr_i[11]
port 536 nsew
rlabel metal2 s 27595 -480 27651 240 4 wbs_adr_i[12]
port 537 nsew
rlabel metal2 s 29389 -480 29445 240 4 wbs_adr_i[13]
port 538 nsew
rlabel metal2 s 31183 -480 31239 240 4 wbs_adr_i[14]
port 539 nsew
rlabel metal2 s 32977 -480 33033 240 4 wbs_adr_i[15]
port 540 nsew
rlabel metal2 s 34725 -480 34781 240 4 wbs_adr_i[16]
port 541 nsew
rlabel metal2 s 36519 -480 36575 240 4 wbs_adr_i[17]
port 542 nsew
rlabel metal2 s 38313 -480 38369 240 4 wbs_adr_i[18]
port 543 nsew
rlabel metal2 s 40107 -480 40163 240 4 wbs_adr_i[19]
port 544 nsew
rlabel metal2 s 6205 -480 6261 240 4 wbs_adr_i[1]
port 545 nsew
rlabel metal2 s 41901 -480 41957 240 4 wbs_adr_i[20]
port 546 nsew
rlabel metal2 s 43649 -480 43705 240 4 wbs_adr_i[21]
port 547 nsew
rlabel metal2 s 45443 -480 45499 240 4 wbs_adr_i[22]
port 548 nsew
rlabel metal2 s 47237 -480 47293 240 4 wbs_adr_i[23]
port 549 nsew
rlabel metal2 s 49031 -480 49087 240 4 wbs_adr_i[24]
port 550 nsew
rlabel metal2 s 50779 -480 50835 240 4 wbs_adr_i[25]
port 551 nsew
rlabel metal2 s 52573 -480 52629 240 4 wbs_adr_i[26]
port 552 nsew
rlabel metal2 s 54367 -480 54423 240 4 wbs_adr_i[27]
port 553 nsew
rlabel metal2 s 56161 -480 56217 240 4 wbs_adr_i[28]
port 554 nsew
rlabel metal2 s 57955 -480 58011 240 4 wbs_adr_i[29]
port 555 nsew
rlabel metal2 s 8597 -480 8653 240 4 wbs_adr_i[2]
port 556 nsew
rlabel metal2 s 59703 -480 59759 240 4 wbs_adr_i[30]
port 557 nsew
rlabel metal2 s 61497 -480 61553 240 4 wbs_adr_i[31]
port 558 nsew
rlabel metal2 s 10943 -480 10999 240 4 wbs_adr_i[3]
port 559 nsew
rlabel metal2 s 13335 -480 13391 240 4 wbs_adr_i[4]
port 560 nsew
rlabel metal2 s 15129 -480 15185 240 4 wbs_adr_i[5]
port 561 nsew
rlabel metal2 s 16923 -480 16979 240 4 wbs_adr_i[6]
port 562 nsew
rlabel metal2 s 18671 -480 18727 240 4 wbs_adr_i[7]
port 563 nsew
rlabel metal2 s 20465 -480 20521 240 4 wbs_adr_i[8]
port 564 nsew
rlabel metal2 s 22259 -480 22315 240 4 wbs_adr_i[9]
port 565 nsew
rlabel metal2 s 2019 -480 2075 240 4 wbs_cyc_i
port 566 nsew
rlabel metal2 s 4411 -480 4467 240 4 wbs_dat_i[0]
port 567 nsew
rlabel metal2 s 24651 -480 24707 240 4 wbs_dat_i[10]
port 568 nsew
rlabel metal2 s 26399 -480 26455 240 4 wbs_dat_i[11]
port 569 nsew
rlabel metal2 s 28193 -480 28249 240 4 wbs_dat_i[12]
port 570 nsew
rlabel metal2 s 29987 -480 30043 240 4 wbs_dat_i[13]
port 571 nsew
rlabel metal2 s 31781 -480 31837 240 4 wbs_dat_i[14]
port 572 nsew
rlabel metal2 s 33575 -480 33631 240 4 wbs_dat_i[15]
port 573 nsew
rlabel metal2 s 35323 -480 35379 240 4 wbs_dat_i[16]
port 574 nsew
rlabel metal2 s 37117 -480 37173 240 4 wbs_dat_i[17]
port 575 nsew
rlabel metal2 s 38911 -480 38967 240 4 wbs_dat_i[18]
port 576 nsew
rlabel metal2 s 40705 -480 40761 240 4 wbs_dat_i[19]
port 577 nsew
rlabel metal2 s 6803 -480 6859 240 4 wbs_dat_i[1]
port 578 nsew
rlabel metal2 s 42453 -480 42509 240 4 wbs_dat_i[20]
port 579 nsew
rlabel metal2 s 44247 -480 44303 240 4 wbs_dat_i[21]
port 580 nsew
rlabel metal2 s 46041 -480 46097 240 4 wbs_dat_i[22]
port 581 nsew
rlabel metal2 s 47835 -480 47891 240 4 wbs_dat_i[23]
port 582 nsew
rlabel metal2 s 49629 -480 49685 240 4 wbs_dat_i[24]
port 583 nsew
rlabel metal2 s 51377 -480 51433 240 4 wbs_dat_i[25]
port 584 nsew
rlabel metal2 s 53171 -480 53227 240 4 wbs_dat_i[26]
port 585 nsew
rlabel metal2 s 54965 -480 55021 240 4 wbs_dat_i[27]
port 586 nsew
rlabel metal2 s 56759 -480 56815 240 4 wbs_dat_i[28]
port 587 nsew
rlabel metal2 s 58553 -480 58609 240 4 wbs_dat_i[29]
port 588 nsew
rlabel metal2 s 9149 -480 9205 240 4 wbs_dat_i[2]
port 589 nsew
rlabel metal2 s 60301 -480 60357 240 4 wbs_dat_i[30]
port 590 nsew
rlabel metal2 s 62095 -480 62151 240 4 wbs_dat_i[31]
port 591 nsew
rlabel metal2 s 11541 -480 11597 240 4 wbs_dat_i[3]
port 592 nsew
rlabel metal2 s 13933 -480 13989 240 4 wbs_dat_i[4]
port 593 nsew
rlabel metal2 s 15727 -480 15783 240 4 wbs_dat_i[5]
port 594 nsew
rlabel metal2 s 17475 -480 17531 240 4 wbs_dat_i[6]
port 595 nsew
rlabel metal2 s 19269 -480 19325 240 4 wbs_dat_i[7]
port 596 nsew
rlabel metal2 s 21063 -480 21119 240 4 wbs_dat_i[8]
port 597 nsew
rlabel metal2 s 22857 -480 22913 240 4 wbs_dat_i[9]
port 598 nsew
rlabel metal2 s 5009 -480 5065 240 4 wbs_dat_o[0]
port 599 nsew
rlabel metal2 s 25249 -480 25305 240 4 wbs_dat_o[10]
port 600 nsew
rlabel metal2 s 26997 -480 27053 240 4 wbs_dat_o[11]
port 601 nsew
rlabel metal2 s 28791 -480 28847 240 4 wbs_dat_o[12]
port 602 nsew
rlabel metal2 s 30585 -480 30641 240 4 wbs_dat_o[13]
port 603 nsew
rlabel metal2 s 32379 -480 32435 240 4 wbs_dat_o[14]
port 604 nsew
rlabel metal2 s 34127 -480 34183 240 4 wbs_dat_o[15]
port 605 nsew
rlabel metal2 s 35921 -480 35977 240 4 wbs_dat_o[16]
port 606 nsew
rlabel metal2 s 37715 -480 37771 240 4 wbs_dat_o[17]
port 607 nsew
rlabel metal2 s 39509 -480 39565 240 4 wbs_dat_o[18]
port 608 nsew
rlabel metal2 s 41303 -480 41359 240 4 wbs_dat_o[19]
port 609 nsew
rlabel metal2 s 7401 -480 7457 240 4 wbs_dat_o[1]
port 610 nsew
rlabel metal2 s 43051 -480 43107 240 4 wbs_dat_o[20]
port 611 nsew
rlabel metal2 s 44845 -480 44901 240 4 wbs_dat_o[21]
port 612 nsew
rlabel metal2 s 46639 -480 46695 240 4 wbs_dat_o[22]
port 613 nsew
rlabel metal2 s 48433 -480 48489 240 4 wbs_dat_o[23]
port 614 nsew
rlabel metal2 s 50227 -480 50283 240 4 wbs_dat_o[24]
port 615 nsew
rlabel metal2 s 51975 -480 52031 240 4 wbs_dat_o[25]
port 616 nsew
rlabel metal2 s 53769 -480 53825 240 4 wbs_dat_o[26]
port 617 nsew
rlabel metal2 s 55563 -480 55619 240 4 wbs_dat_o[27]
port 618 nsew
rlabel metal2 s 57357 -480 57413 240 4 wbs_dat_o[28]
port 619 nsew
rlabel metal2 s 59105 -480 59161 240 4 wbs_dat_o[29]
port 620 nsew
rlabel metal2 s 9747 -480 9803 240 4 wbs_dat_o[2]
port 621 nsew
rlabel metal2 s 60899 -480 60955 240 4 wbs_dat_o[30]
port 622 nsew
rlabel metal2 s 62693 -480 62749 240 4 wbs_dat_o[31]
port 623 nsew
rlabel metal2 s 12139 -480 12195 240 4 wbs_dat_o[3]
port 624 nsew
rlabel metal2 s 14531 -480 14587 240 4 wbs_dat_o[4]
port 625 nsew
rlabel metal2 s 16325 -480 16381 240 4 wbs_dat_o[5]
port 626 nsew
rlabel metal2 s 18073 -480 18129 240 4 wbs_dat_o[6]
port 627 nsew
rlabel metal2 s 19867 -480 19923 240 4 wbs_dat_o[7]
port 628 nsew
rlabel metal2 s 21661 -480 21717 240 4 wbs_dat_o[8]
port 629 nsew
rlabel metal2 s 23455 -480 23511 240 4 wbs_dat_o[9]
port 630 nsew
rlabel metal2 s 5607 -480 5663 240 4 wbs_sel_i[0]
port 631 nsew
rlabel metal2 s 7999 -480 8055 240 4 wbs_sel_i[1]
port 632 nsew
rlabel metal2 s 10345 -480 10401 240 4 wbs_sel_i[2]
port 633 nsew
rlabel metal2 s 12737 -480 12793 240 4 wbs_sel_i[3]
port 634 nsew
rlabel metal2 s 2617 -480 2673 240 4 wbs_stb_i
port 635 nsew
rlabel metal2 s 3215 -480 3271 240 4 wbs_we_i
port 636 nsew
rlabel metal5 s -998 -462 292960 -162 4 vccd1
port 637 nsew
rlabel metal5 s -1458 -922 293420 -622 4 vssd1
port 638 nsew
rlabel metal5 s -1918 -1382 293880 -1082 4 vccd2
port 639 nsew
rlabel metal5 s -2378 -1842 294340 -1542 4 vssd2
port 640 nsew
rlabel metal5 s -2838 -2302 294800 -2002 4 vdda1
port 641 nsew
rlabel metal5 s -3298 -2762 295260 -2462 4 vssa1
port 642 nsew
rlabel metal5 s -3758 -3222 295720 -2922 4 vdda2
port 643 nsew
rlabel metal5 s -4218 -3682 296180 -3382 4 vssa2
port 644 nsew
<< properties >>
string FIXED_BBOX 0 0 292000 352000
string GDS_FILE /project/openlane/user_project_wrapper_empty/runs/user_project_wrapper_empty/results/magic/user_project_wrapper.gds
string GDS_END 306838
string GDS_START 130
<< end >>
