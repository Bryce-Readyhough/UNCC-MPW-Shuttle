magic
tech sky130A
timestamp 1606420262
<< metal2 >>
rect 4793 269760 4821 270000
rect 14407 269760 14435 270000
rect 24067 269760 24095 270000
rect 33681 269760 33709 270000
rect 43341 269760 43369 270000
rect 53001 269760 53029 270000
rect 62615 269760 62643 270000
rect 72275 269760 72303 270000
rect 81935 269760 81963 270000
rect 91549 269760 91577 270000
rect 101209 269760 101237 270000
rect 110869 269760 110897 270000
rect 120483 269760 120511 270000
rect 130143 269760 130171 270000
rect 139803 269760 139831 270000
rect 149417 269760 149445 270000
rect 159077 269760 159105 270000
rect 168691 269760 168719 270000
rect 178351 269760 178379 270000
rect 188011 269760 188039 270000
rect 197625 269760 197653 270000
rect 207285 269760 207313 270000
rect 216945 269760 216973 270000
rect 226559 269760 226587 270000
rect 236219 269760 236247 270000
rect 245879 269760 245907 270000
rect 255493 269760 255521 270000
rect 265153 269760 265181 270000
rect 239 0 267 240
rect 745 0 773 240
rect 1297 0 1325 240
rect 1849 0 1877 240
rect 2401 0 2429 240
rect 2953 0 2981 240
rect 3505 0 3533 240
rect 4057 0 4085 240
rect 4609 0 4637 240
rect 5161 0 5189 240
rect 5713 0 5741 240
rect 6265 0 6293 240
rect 6817 0 6845 240
rect 7369 0 7397 240
rect 7921 0 7949 240
rect 8473 0 8501 240
rect 9025 0 9053 240
rect 9577 0 9605 240
rect 10129 0 10157 240
rect 10681 0 10709 240
rect 11233 0 11261 240
rect 11785 0 11813 240
rect 12337 0 12365 240
rect 12843 0 12871 240
rect 13395 0 13423 240
rect 13947 0 13975 240
rect 14499 0 14527 240
rect 15051 0 15079 240
rect 15603 0 15631 240
rect 16155 0 16183 240
rect 16707 0 16735 240
rect 17259 0 17287 240
rect 17811 0 17839 240
rect 18363 0 18391 240
rect 18915 0 18943 240
rect 19467 0 19495 240
rect 20019 0 20047 240
rect 20571 0 20599 240
rect 21123 0 21151 240
rect 21675 0 21703 240
rect 22227 0 22255 240
rect 22779 0 22807 240
rect 23331 0 23359 240
rect 23883 0 23911 240
rect 24435 0 24463 240
rect 24941 0 24969 240
rect 25493 0 25521 240
rect 26045 0 26073 240
rect 26597 0 26625 240
rect 27149 0 27177 240
rect 27701 0 27729 240
rect 28253 0 28281 240
rect 28805 0 28833 240
rect 29357 0 29385 240
rect 29909 0 29937 240
rect 30461 0 30489 240
rect 31013 0 31041 240
rect 31565 0 31593 240
rect 32117 0 32145 240
rect 32669 0 32697 240
rect 33221 0 33249 240
rect 33773 0 33801 240
rect 34325 0 34353 240
rect 34877 0 34905 240
rect 35429 0 35457 240
rect 35981 0 36009 240
rect 36533 0 36561 240
rect 37039 0 37067 240
rect 37591 0 37619 240
rect 38143 0 38171 240
rect 38695 0 38723 240
rect 39247 0 39275 240
rect 39799 0 39827 240
rect 40351 0 40379 240
rect 40903 0 40931 240
rect 41455 0 41483 240
rect 42007 0 42035 240
rect 42559 0 42587 240
rect 43111 0 43139 240
rect 43663 0 43691 240
rect 44215 0 44243 240
rect 44767 0 44795 240
rect 45319 0 45347 240
rect 45871 0 45899 240
rect 46423 0 46451 240
rect 46975 0 47003 240
rect 47527 0 47555 240
rect 48079 0 48107 240
rect 48631 0 48659 240
rect 49183 0 49211 240
rect 49689 0 49717 240
rect 50241 0 50269 240
rect 50793 0 50821 240
rect 51345 0 51373 240
rect 51897 0 51925 240
rect 52449 0 52477 240
rect 53001 0 53029 240
rect 53553 0 53581 240
rect 54105 0 54133 240
rect 54657 0 54685 240
rect 55209 0 55237 240
rect 55761 0 55789 240
rect 56313 0 56341 240
rect 56865 0 56893 240
rect 57417 0 57445 240
rect 57969 0 57997 240
rect 58521 0 58549 240
rect 59073 0 59101 240
rect 59625 0 59653 240
rect 60177 0 60205 240
rect 60729 0 60757 240
rect 61281 0 61309 240
rect 61787 0 61815 240
rect 62339 0 62367 240
rect 62891 0 62919 240
rect 63443 0 63471 240
rect 63995 0 64023 240
rect 64547 0 64575 240
rect 65099 0 65127 240
rect 65651 0 65679 240
rect 66203 0 66231 240
rect 66755 0 66783 240
rect 67307 0 67335 240
rect 67859 0 67887 240
rect 68411 0 68439 240
rect 68963 0 68991 240
rect 69515 0 69543 240
rect 70067 0 70095 240
rect 70619 0 70647 240
rect 71171 0 71199 240
rect 71723 0 71751 240
rect 72275 0 72303 240
rect 72827 0 72855 240
rect 73379 0 73407 240
rect 73885 0 73913 240
rect 74437 0 74465 240
rect 74989 0 75017 240
rect 75541 0 75569 240
rect 76093 0 76121 240
rect 76645 0 76673 240
rect 77197 0 77225 240
rect 77749 0 77777 240
rect 78301 0 78329 240
rect 78853 0 78881 240
rect 79405 0 79433 240
rect 79957 0 79985 240
rect 80509 0 80537 240
rect 81061 0 81089 240
rect 81613 0 81641 240
rect 82165 0 82193 240
rect 82717 0 82745 240
rect 83269 0 83297 240
rect 83821 0 83849 240
rect 84373 0 84401 240
rect 84925 0 84953 240
rect 85477 0 85505 240
rect 86029 0 86057 240
rect 86535 0 86563 240
rect 87087 0 87115 240
rect 87639 0 87667 240
rect 88191 0 88219 240
rect 88743 0 88771 240
rect 89295 0 89323 240
rect 89847 0 89875 240
rect 90399 0 90427 240
rect 90951 0 90979 240
rect 91503 0 91531 240
rect 92055 0 92083 240
rect 92607 0 92635 240
rect 93159 0 93187 240
rect 93711 0 93739 240
rect 94263 0 94291 240
rect 94815 0 94843 240
rect 95367 0 95395 240
rect 95919 0 95947 240
rect 96471 0 96499 240
rect 97023 0 97051 240
rect 97575 0 97603 240
rect 98127 0 98155 240
rect 98633 0 98661 240
rect 99185 0 99213 240
rect 99737 0 99765 240
rect 100289 0 100317 240
rect 100841 0 100869 240
rect 101393 0 101421 240
rect 101945 0 101973 240
rect 102497 0 102525 240
rect 103049 0 103077 240
rect 103601 0 103629 240
rect 104153 0 104181 240
rect 104705 0 104733 240
rect 105257 0 105285 240
rect 105809 0 105837 240
rect 106361 0 106389 240
rect 106913 0 106941 240
rect 107465 0 107493 240
rect 108017 0 108045 240
rect 108569 0 108597 240
rect 109121 0 109149 240
rect 109673 0 109701 240
rect 110225 0 110253 240
rect 110731 0 110759 240
rect 111283 0 111311 240
rect 111835 0 111863 240
rect 112387 0 112415 240
rect 112939 0 112967 240
rect 113491 0 113519 240
rect 114043 0 114071 240
rect 114595 0 114623 240
rect 115147 0 115175 240
rect 115699 0 115727 240
rect 116251 0 116279 240
rect 116803 0 116831 240
rect 117355 0 117383 240
rect 117907 0 117935 240
rect 118459 0 118487 240
rect 119011 0 119039 240
rect 119563 0 119591 240
rect 120115 0 120143 240
rect 120667 0 120695 240
rect 121219 0 121247 240
rect 121771 0 121799 240
rect 122323 0 122351 240
rect 122875 0 122903 240
rect 123381 0 123409 240
rect 123933 0 123961 240
rect 124485 0 124513 240
rect 125037 0 125065 240
rect 125589 0 125617 240
rect 126141 0 126169 240
rect 126693 0 126721 240
rect 127245 0 127273 240
rect 127797 0 127825 240
rect 128349 0 128377 240
rect 128901 0 128929 240
rect 129453 0 129481 240
rect 130005 0 130033 240
rect 130557 0 130585 240
rect 131109 0 131137 240
rect 131661 0 131689 240
rect 132213 0 132241 240
rect 132765 0 132793 240
rect 133317 0 133345 240
rect 133869 0 133897 240
rect 134421 0 134449 240
rect 134973 0 135001 240
rect 135479 0 135507 240
rect 136031 0 136059 240
rect 136583 0 136611 240
rect 137135 0 137163 240
rect 137687 0 137715 240
rect 138239 0 138267 240
rect 138791 0 138819 240
rect 139343 0 139371 240
rect 139895 0 139923 240
rect 140447 0 140475 240
rect 140999 0 141027 240
rect 141551 0 141579 240
rect 142103 0 142131 240
rect 142655 0 142683 240
rect 143207 0 143235 240
rect 143759 0 143787 240
rect 144311 0 144339 240
rect 144863 0 144891 240
rect 145415 0 145443 240
rect 145967 0 145995 240
rect 146519 0 146547 240
rect 147071 0 147099 240
rect 147577 0 147605 240
rect 148129 0 148157 240
rect 148681 0 148709 240
rect 149233 0 149261 240
rect 149785 0 149813 240
rect 150337 0 150365 240
rect 150889 0 150917 240
rect 151441 0 151469 240
rect 151993 0 152021 240
rect 152545 0 152573 240
rect 153097 0 153125 240
rect 153649 0 153677 240
rect 154201 0 154229 240
rect 154753 0 154781 240
rect 155305 0 155333 240
rect 155857 0 155885 240
rect 156409 0 156437 240
rect 156961 0 156989 240
rect 157513 0 157541 240
rect 158065 0 158093 240
rect 158617 0 158645 240
rect 159169 0 159197 240
rect 159721 0 159749 240
rect 160227 0 160255 240
rect 160779 0 160807 240
rect 161331 0 161359 240
rect 161883 0 161911 240
rect 162435 0 162463 240
rect 162987 0 163015 240
rect 163539 0 163567 240
rect 164091 0 164119 240
rect 164643 0 164671 240
rect 165195 0 165223 240
rect 165747 0 165775 240
rect 166299 0 166327 240
rect 166851 0 166879 240
rect 167403 0 167431 240
rect 167955 0 167983 240
rect 168507 0 168535 240
rect 169059 0 169087 240
rect 169611 0 169639 240
rect 170163 0 170191 240
rect 170715 0 170743 240
rect 171267 0 171295 240
rect 171819 0 171847 240
rect 172325 0 172353 240
rect 172877 0 172905 240
rect 173429 0 173457 240
rect 173981 0 174009 240
rect 174533 0 174561 240
rect 175085 0 175113 240
rect 175637 0 175665 240
rect 176189 0 176217 240
rect 176741 0 176769 240
rect 177293 0 177321 240
rect 177845 0 177873 240
rect 178397 0 178425 240
rect 178949 0 178977 240
rect 179501 0 179529 240
rect 180053 0 180081 240
rect 180605 0 180633 240
rect 181157 0 181185 240
rect 181709 0 181737 240
rect 182261 0 182289 240
rect 182813 0 182841 240
rect 183365 0 183393 240
rect 183917 0 183945 240
rect 184423 0 184451 240
rect 184975 0 185003 240
rect 185527 0 185555 240
rect 186079 0 186107 240
rect 186631 0 186659 240
rect 187183 0 187211 240
rect 187735 0 187763 240
rect 188287 0 188315 240
rect 188839 0 188867 240
rect 189391 0 189419 240
rect 189943 0 189971 240
rect 190495 0 190523 240
rect 191047 0 191075 240
rect 191599 0 191627 240
rect 192151 0 192179 240
rect 192703 0 192731 240
rect 193255 0 193283 240
rect 193807 0 193835 240
rect 194359 0 194387 240
rect 194911 0 194939 240
rect 195463 0 195491 240
rect 196015 0 196043 240
rect 196567 0 196595 240
rect 197073 0 197101 240
rect 197625 0 197653 240
rect 198177 0 198205 240
rect 198729 0 198757 240
rect 199281 0 199309 240
rect 199833 0 199861 240
rect 200385 0 200413 240
rect 200937 0 200965 240
rect 201489 0 201517 240
rect 202041 0 202069 240
rect 202593 0 202621 240
rect 203145 0 203173 240
rect 203697 0 203725 240
rect 204249 0 204277 240
rect 204801 0 204829 240
rect 205353 0 205381 240
rect 205905 0 205933 240
rect 206457 0 206485 240
rect 207009 0 207037 240
rect 207561 0 207589 240
rect 208113 0 208141 240
rect 208665 0 208693 240
rect 209171 0 209199 240
rect 209723 0 209751 240
rect 210275 0 210303 240
rect 210827 0 210855 240
rect 211379 0 211407 240
rect 211931 0 211959 240
rect 212483 0 212511 240
rect 213035 0 213063 240
rect 213587 0 213615 240
rect 214139 0 214167 240
rect 214691 0 214719 240
rect 215243 0 215271 240
rect 215795 0 215823 240
rect 216347 0 216375 240
rect 216899 0 216927 240
rect 217451 0 217479 240
rect 218003 0 218031 240
rect 218555 0 218583 240
rect 219107 0 219135 240
rect 219659 0 219687 240
rect 220211 0 220239 240
rect 220763 0 220791 240
rect 221269 0 221297 240
rect 221821 0 221849 240
rect 222373 0 222401 240
rect 222925 0 222953 240
rect 223477 0 223505 240
rect 224029 0 224057 240
rect 224581 0 224609 240
rect 225133 0 225161 240
rect 225685 0 225713 240
rect 226237 0 226265 240
rect 226789 0 226817 240
rect 227341 0 227369 240
rect 227893 0 227921 240
rect 228445 0 228473 240
rect 228997 0 229025 240
rect 229549 0 229577 240
rect 230101 0 230129 240
rect 230653 0 230681 240
rect 231205 0 231233 240
rect 231757 0 231785 240
rect 232309 0 232337 240
rect 232861 0 232889 240
rect 233413 0 233441 240
rect 233919 0 233947 240
rect 234471 0 234499 240
rect 235023 0 235051 240
rect 235575 0 235603 240
rect 236127 0 236155 240
rect 236679 0 236707 240
rect 237231 0 237259 240
rect 237783 0 237811 240
rect 238335 0 238363 240
rect 238887 0 238915 240
rect 239439 0 239467 240
rect 239991 0 240019 240
rect 240543 0 240571 240
rect 241095 0 241123 240
rect 241647 0 241675 240
rect 242199 0 242227 240
rect 242751 0 242779 240
rect 243303 0 243331 240
rect 243855 0 243883 240
rect 244407 0 244435 240
rect 244959 0 244987 240
rect 245511 0 245539 240
rect 246017 0 246045 240
rect 246569 0 246597 240
rect 247121 0 247149 240
rect 247673 0 247701 240
rect 248225 0 248253 240
rect 248777 0 248805 240
rect 249329 0 249357 240
rect 249881 0 249909 240
rect 250433 0 250461 240
rect 250985 0 251013 240
rect 251537 0 251565 240
rect 252089 0 252117 240
rect 252641 0 252669 240
rect 253193 0 253221 240
rect 253745 0 253773 240
rect 254297 0 254325 240
rect 254849 0 254877 240
rect 255401 0 255429 240
rect 255953 0 255981 240
rect 256505 0 256533 240
rect 257057 0 257085 240
rect 257609 0 257637 240
rect 258115 0 258143 240
rect 258667 0 258695 240
rect 259219 0 259247 240
rect 259771 0 259799 240
rect 260323 0 260351 240
rect 260875 0 260903 240
rect 261427 0 261455 240
rect 261979 0 262007 240
rect 262531 0 262559 240
rect 263083 0 263111 240
rect 263635 0 263663 240
rect 264187 0 264215 240
rect 264739 0 264767 240
rect 265291 0 265319 240
rect 265843 0 265871 240
rect 266395 0 266423 240
rect 266947 0 266975 240
rect 267499 0 267527 240
rect 268051 0 268079 240
rect 268603 0 268631 240
rect 269155 0 269183 240
rect 269707 0 269735 240
<< metal3 >>
rect 269760 267176 270000 267236
rect 0 267040 240 267100
rect 269760 261532 270000 261592
rect 0 261192 240 261252
rect 269760 255888 270000 255948
rect 0 255344 240 255404
rect 269760 250312 270000 250372
rect 0 249428 240 249488
rect 269760 244668 270000 244728
rect 0 243580 240 243640
rect 269760 239024 270000 239084
rect 0 237732 240 237792
rect 269760 233380 270000 233440
rect 0 231816 240 231876
rect 269760 227804 270000 227864
rect 0 225968 240 226028
rect 269760 222160 270000 222220
rect 0 220120 240 220180
rect 269760 216516 270000 216576
rect 0 214204 240 214264
rect 269760 210872 270000 210932
rect 0 208356 240 208416
rect 269760 205296 270000 205356
rect 0 202508 240 202568
rect 269760 199652 270000 199712
rect 0 196592 240 196652
rect 269760 194008 270000 194068
rect 0 190744 240 190804
rect 269760 188432 270000 188492
rect 0 184896 240 184956
rect 269760 182788 270000 182848
rect 0 178980 240 179040
rect 269760 177144 270000 177204
rect 0 173132 240 173192
rect 269760 171500 270000 171560
rect 0 167284 240 167344
rect 269760 165924 270000 165984
rect 0 161368 240 161428
rect 269760 160280 270000 160340
rect 0 155520 240 155580
rect 269760 154636 270000 154696
rect 0 149672 240 149732
rect 269760 148992 270000 149052
rect 0 143756 240 143816
rect 269760 143416 270000 143476
rect 0 137908 240 137968
rect 269760 137772 270000 137832
rect 269760 132128 270000 132188
rect 0 132060 240 132120
rect 269760 126552 270000 126612
rect 0 126144 240 126204
rect 269760 120908 270000 120968
rect 0 120296 240 120356
rect 269760 115264 270000 115324
rect 0 114448 240 114508
rect 269760 109620 270000 109680
rect 0 108532 240 108592
rect 269760 104044 270000 104104
rect 0 102684 240 102744
rect 269760 98400 270000 98460
rect 0 96836 240 96896
rect 269760 92756 270000 92816
rect 0 90920 240 90980
rect 269760 87112 270000 87172
rect 0 85072 240 85132
rect 269760 81536 270000 81596
rect 0 79224 240 79284
rect 269760 75892 270000 75952
rect 0 73308 240 73368
rect 269760 70248 270000 70308
rect 0 67460 240 67520
rect 269760 64672 270000 64732
rect 0 61612 240 61672
rect 269760 59028 270000 59088
rect 0 55696 240 55756
rect 269760 53384 270000 53444
rect 0 49848 240 49908
rect 269760 47740 270000 47800
rect 0 44000 240 44060
rect 269760 42164 270000 42224
rect 0 38084 240 38144
rect 269760 36520 270000 36580
rect 0 32236 240 32296
rect 269760 30876 270000 30936
rect 0 26388 240 26448
rect 269760 25232 270000 25292
rect 0 20472 240 20532
rect 269760 19656 270000 19716
rect 0 14624 240 14684
rect 269760 14012 270000 14072
rect 0 8776 240 8836
rect 269760 8368 270000 8428
rect 0 2928 240 2988
rect 269760 2792 270000 2852
use chip-2  chip-2_0 ~/UNCCCaravel/UNCC-MPW-Shuttle/mag/tinysky
timestamp 1606345435
transform 1 0 150722 0 1 76312
box -12242 -4023 9920 9117
<< labels >>
rlabel metal3 s 269760 2792 270000 2852 6 io_in[0]
port 0 nsew default input
rlabel metal3 s 269760 182788 270000 182848 6 io_in[10]
port 1 nsew default input
rlabel metal3 s 269760 199652 270000 199712 6 io_in[11]
port 2 nsew default input
rlabel metal3 s 269760 216516 270000 216576 6 io_in[12]
port 3 nsew default input
rlabel metal3 s 269760 233380 270000 233440 6 io_in[13]
port 4 nsew default input
rlabel metal3 s 269760 255888 270000 255948 6 io_in[14]
port 5 nsew default input
rlabel metal2 s 265153 269760 265181 270000 6 io_in[15]
port 6 nsew default input
rlabel metal2 s 226559 269760 226587 270000 6 io_in[16]
port 7 nsew default input
rlabel metal2 s 197625 269760 197653 270000 6 io_in[17]
port 8 nsew default input
rlabel metal2 s 168691 269760 168719 270000 6 io_in[18]
port 9 nsew default input
rlabel metal2 s 139803 269760 139831 270000 6 io_in[19]
port 10 nsew default input
rlabel metal3 s 269760 19656 270000 19716 6 io_in[1]
port 11 nsew default input
rlabel metal2 s 110869 269760 110897 270000 6 io_in[20]
port 12 nsew default input
rlabel metal2 s 81935 269760 81963 270000 6 io_in[21]
port 13 nsew default input
rlabel metal2 s 53001 269760 53029 270000 6 io_in[22]
port 14 nsew default input
rlabel metal2 s 24067 269760 24095 270000 6 io_in[23]
port 15 nsew default input
rlabel metal3 s 0 267040 240 267100 6 io_in[24]
port 16 nsew default input
rlabel metal3 s 0 237732 240 237792 6 io_in[25]
port 17 nsew default input
rlabel metal3 s 0 220120 240 220180 6 io_in[26]
port 18 nsew default input
rlabel metal3 s 0 202508 240 202568 6 io_in[27]
port 19 nsew default input
rlabel metal3 s 0 184896 240 184956 6 io_in[28]
port 20 nsew default input
rlabel metal3 s 0 167284 240 167344 6 io_in[29]
port 21 nsew default input
rlabel metal3 s 269760 36520 270000 36580 6 io_in[2]
port 22 nsew default input
rlabel metal3 s 0 149672 240 149732 6 io_in[30]
port 23 nsew default input
rlabel metal3 s 0 132060 240 132120 6 io_in[31]
port 24 nsew default input
rlabel metal3 s 0 102684 240 102744 6 io_in[32]
port 25 nsew default input
rlabel metal3 s 0 85072 240 85132 6 io_in[33]
port 26 nsew default input
rlabel metal3 s 0 67460 240 67520 6 io_in[34]
port 27 nsew default input
rlabel metal3 s 0 49848 240 49908 6 io_in[35]
port 28 nsew default input
rlabel metal3 s 0 32236 240 32296 6 io_in[36]
port 29 nsew default input
rlabel metal3 s 0 14624 240 14684 6 io_in[37]
port 30 nsew default input
rlabel metal3 s 269760 53384 270000 53444 6 io_in[3]
port 31 nsew default input
rlabel metal3 s 269760 70248 270000 70308 6 io_in[4]
port 32 nsew default input
rlabel metal3 s 269760 87112 270000 87172 6 io_in[5]
port 33 nsew default input
rlabel metal3 s 269760 104044 270000 104104 6 io_in[6]
port 34 nsew default input
rlabel metal3 s 269760 132128 270000 132188 6 io_in[7]
port 35 nsew default input
rlabel metal3 s 269760 148992 270000 149052 6 io_in[8]
port 36 nsew default input
rlabel metal3 s 269760 165924 270000 165984 6 io_in[9]
port 37 nsew default input
rlabel metal3 s 269760 14012 270000 14072 6 io_oeb[0]
port 38 nsew default tristate
rlabel metal3 s 269760 194008 270000 194068 6 io_oeb[10]
port 39 nsew default tristate
rlabel metal3 s 269760 210872 270000 210932 6 io_oeb[11]
port 40 nsew default tristate
rlabel metal3 s 269760 227804 270000 227864 6 io_oeb[12]
port 41 nsew default tristate
rlabel metal3 s 269760 244668 270000 244728 6 io_oeb[13]
port 42 nsew default tristate
rlabel metal3 s 269760 267176 270000 267236 6 io_oeb[14]
port 43 nsew default tristate
rlabel metal2 s 245879 269760 245907 270000 6 io_oeb[15]
port 44 nsew default tristate
rlabel metal2 s 207285 269760 207313 270000 6 io_oeb[16]
port 45 nsew default tristate
rlabel metal2 s 178351 269760 178379 270000 6 io_oeb[17]
port 46 nsew default tristate
rlabel metal2 s 149417 269760 149445 270000 6 io_oeb[18]
port 47 nsew default tristate
rlabel metal2 s 120483 269760 120511 270000 6 io_oeb[19]
port 48 nsew default tristate
rlabel metal3 s 269760 30876 270000 30936 6 io_oeb[1]
port 49 nsew default tristate
rlabel metal2 s 91549 269760 91577 270000 6 io_oeb[20]
port 50 nsew default tristate
rlabel metal2 s 62615 269760 62643 270000 6 io_oeb[21]
port 51 nsew default tristate
rlabel metal2 s 33681 269760 33709 270000 6 io_oeb[22]
port 52 nsew default tristate
rlabel metal2 s 4793 269760 4821 270000 6 io_oeb[23]
port 53 nsew default tristate
rlabel metal3 s 0 255344 240 255404 6 io_oeb[24]
port 54 nsew default tristate
rlabel metal3 s 0 225968 240 226028 6 io_oeb[25]
port 55 nsew default tristate
rlabel metal3 s 0 208356 240 208416 6 io_oeb[26]
port 56 nsew default tristate
rlabel metal3 s 0 190744 240 190804 6 io_oeb[27]
port 57 nsew default tristate
rlabel metal3 s 0 173132 240 173192 6 io_oeb[28]
port 58 nsew default tristate
rlabel metal3 s 0 155520 240 155580 6 io_oeb[29]
port 59 nsew default tristate
rlabel metal3 s 269760 47740 270000 47800 6 io_oeb[2]
port 60 nsew default tristate
rlabel metal3 s 0 137908 240 137968 6 io_oeb[30]
port 61 nsew default tristate
rlabel metal3 s 0 120296 240 120356 6 io_oeb[31]
port 62 nsew default tristate
rlabel metal3 s 0 90920 240 90980 6 io_oeb[32]
port 63 nsew default tristate
rlabel metal3 s 0 73308 240 73368 6 io_oeb[33]
port 64 nsew default tristate
rlabel metal3 s 0 55696 240 55756 6 io_oeb[34]
port 65 nsew default tristate
rlabel metal3 s 0 38084 240 38144 6 io_oeb[35]
port 66 nsew default tristate
rlabel metal3 s 0 20472 240 20532 6 io_oeb[36]
port 67 nsew default tristate
rlabel metal3 s 0 2928 240 2988 6 io_oeb[37]
port 68 nsew default tristate
rlabel metal3 s 269760 64672 270000 64732 6 io_oeb[3]
port 69 nsew default tristate
rlabel metal3 s 269760 81536 270000 81596 6 io_oeb[4]
port 70 nsew default tristate
rlabel metal3 s 269760 98400 270000 98460 6 io_oeb[5]
port 71 nsew default tristate
rlabel metal3 s 269760 115264 270000 115324 6 io_oeb[6]
port 72 nsew default tristate
rlabel metal3 s 269760 143416 270000 143476 6 io_oeb[7]
port 73 nsew default tristate
rlabel metal3 s 269760 160280 270000 160340 6 io_oeb[8]
port 74 nsew default tristate
rlabel metal3 s 269760 177144 270000 177204 6 io_oeb[9]
port 75 nsew default tristate
rlabel metal3 s 269760 8368 270000 8428 6 io_out[0]
port 76 nsew default tristate
rlabel metal3 s 269760 188432 270000 188492 6 io_out[10]
port 77 nsew default tristate
rlabel metal3 s 269760 205296 270000 205356 6 io_out[11]
port 78 nsew default tristate
rlabel metal3 s 269760 222160 270000 222220 6 io_out[12]
port 79 nsew default tristate
rlabel metal3 s 269760 239024 270000 239084 6 io_out[13]
port 80 nsew default tristate
rlabel metal3 s 269760 261532 270000 261592 6 io_out[14]
port 81 nsew default tristate
rlabel metal2 s 255493 269760 255521 270000 6 io_out[15]
port 82 nsew default tristate
rlabel metal2 s 216945 269760 216973 270000 6 io_out[16]
port 83 nsew default tristate
rlabel metal2 s 188011 269760 188039 270000 6 io_out[17]
port 84 nsew default tristate
rlabel metal2 s 159077 269760 159105 270000 6 io_out[18]
port 85 nsew default tristate
rlabel metal2 s 130143 269760 130171 270000 6 io_out[19]
port 86 nsew default tristate
rlabel metal3 s 269760 25232 270000 25292 6 io_out[1]
port 87 nsew default tristate
rlabel metal2 s 101209 269760 101237 270000 6 io_out[20]
port 88 nsew default tristate
rlabel metal2 s 72275 269760 72303 270000 6 io_out[21]
port 89 nsew default tristate
rlabel metal2 s 43341 269760 43369 270000 6 io_out[22]
port 90 nsew default tristate
rlabel metal2 s 14407 269760 14435 270000 6 io_out[23]
port 91 nsew default tristate
rlabel metal3 s 0 261192 240 261252 6 io_out[24]
port 92 nsew default tristate
rlabel metal3 s 0 231816 240 231876 6 io_out[25]
port 93 nsew default tristate
rlabel metal3 s 0 214204 240 214264 6 io_out[26]
port 94 nsew default tristate
rlabel metal3 s 0 196592 240 196652 6 io_out[27]
port 95 nsew default tristate
rlabel metal3 s 0 178980 240 179040 6 io_out[28]
port 96 nsew default tristate
rlabel metal3 s 0 161368 240 161428 6 io_out[29]
port 97 nsew default tristate
rlabel metal3 s 269760 42164 270000 42224 6 io_out[2]
port 98 nsew default tristate
rlabel metal3 s 0 143756 240 143816 6 io_out[30]
port 99 nsew default tristate
rlabel metal3 s 0 126144 240 126204 6 io_out[31]
port 100 nsew default tristate
rlabel metal3 s 0 96836 240 96896 6 io_out[32]
port 101 nsew default tristate
rlabel metal3 s 0 79224 240 79284 6 io_out[33]
port 102 nsew default tristate
rlabel metal3 s 0 61612 240 61672 6 io_out[34]
port 103 nsew default tristate
rlabel metal3 s 0 44000 240 44060 6 io_out[35]
port 104 nsew default tristate
rlabel metal3 s 0 26388 240 26448 6 io_out[36]
port 105 nsew default tristate
rlabel metal3 s 0 8776 240 8836 6 io_out[37]
port 106 nsew default tristate
rlabel metal3 s 269760 59028 270000 59088 6 io_out[3]
port 107 nsew default tristate
rlabel metal3 s 269760 75892 270000 75952 6 io_out[4]
port 108 nsew default tristate
rlabel metal3 s 269760 92756 270000 92816 6 io_out[5]
port 109 nsew default tristate
rlabel metal3 s 269760 109620 270000 109680 6 io_out[6]
port 110 nsew default tristate
rlabel metal3 s 269760 137772 270000 137832 6 io_out[7]
port 111 nsew default tristate
rlabel metal3 s 269760 154636 270000 154696 6 io_out[8]
port 112 nsew default tristate
rlabel metal3 s 269760 171500 270000 171560 6 io_out[9]
port 113 nsew default tristate
rlabel metal2 s 58521 0 58549 240 6 la_data_in[0]
port 114 nsew default input
rlabel metal2 s 223477 0 223505 240 6 la_data_in[100]
port 115 nsew default input
rlabel metal2 s 225133 0 225161 240 6 la_data_in[101]
port 116 nsew default input
rlabel metal2 s 226789 0 226817 240 6 la_data_in[102]
port 117 nsew default input
rlabel metal2 s 228445 0 228473 240 6 la_data_in[103]
port 118 nsew default input
rlabel metal2 s 230101 0 230129 240 6 la_data_in[104]
port 119 nsew default input
rlabel metal2 s 231757 0 231785 240 6 la_data_in[105]
port 120 nsew default input
rlabel metal2 s 233413 0 233441 240 6 la_data_in[106]
port 121 nsew default input
rlabel metal2 s 235023 0 235051 240 6 la_data_in[107]
port 122 nsew default input
rlabel metal2 s 236679 0 236707 240 6 la_data_in[108]
port 123 nsew default input
rlabel metal2 s 238335 0 238363 240 6 la_data_in[109]
port 124 nsew default input
rlabel metal2 s 74989 0 75017 240 6 la_data_in[10]
port 125 nsew default input
rlabel metal2 s 239991 0 240019 240 6 la_data_in[110]
port 126 nsew default input
rlabel metal2 s 241647 0 241675 240 6 la_data_in[111]
port 127 nsew default input
rlabel metal2 s 243303 0 243331 240 6 la_data_in[112]
port 128 nsew default input
rlabel metal2 s 244959 0 244987 240 6 la_data_in[113]
port 129 nsew default input
rlabel metal2 s 246569 0 246597 240 6 la_data_in[114]
port 130 nsew default input
rlabel metal2 s 248225 0 248253 240 6 la_data_in[115]
port 131 nsew default input
rlabel metal2 s 249881 0 249909 240 6 la_data_in[116]
port 132 nsew default input
rlabel metal2 s 251537 0 251565 240 6 la_data_in[117]
port 133 nsew default input
rlabel metal2 s 253193 0 253221 240 6 la_data_in[118]
port 134 nsew default input
rlabel metal2 s 254849 0 254877 240 6 la_data_in[119]
port 135 nsew default input
rlabel metal2 s 76645 0 76673 240 6 la_data_in[11]
port 136 nsew default input
rlabel metal2 s 256505 0 256533 240 6 la_data_in[120]
port 137 nsew default input
rlabel metal2 s 258115 0 258143 240 6 la_data_in[121]
port 138 nsew default input
rlabel metal2 s 259771 0 259799 240 6 la_data_in[122]
port 139 nsew default input
rlabel metal2 s 261427 0 261455 240 6 la_data_in[123]
port 140 nsew default input
rlabel metal2 s 263083 0 263111 240 6 la_data_in[124]
port 141 nsew default input
rlabel metal2 s 264739 0 264767 240 6 la_data_in[125]
port 142 nsew default input
rlabel metal2 s 266395 0 266423 240 6 la_data_in[126]
port 143 nsew default input
rlabel metal2 s 268051 0 268079 240 6 la_data_in[127]
port 144 nsew default input
rlabel metal2 s 78301 0 78329 240 6 la_data_in[12]
port 145 nsew default input
rlabel metal2 s 79957 0 79985 240 6 la_data_in[13]
port 146 nsew default input
rlabel metal2 s 81613 0 81641 240 6 la_data_in[14]
port 147 nsew default input
rlabel metal2 s 83269 0 83297 240 6 la_data_in[15]
port 148 nsew default input
rlabel metal2 s 84925 0 84953 240 6 la_data_in[16]
port 149 nsew default input
rlabel metal2 s 86535 0 86563 240 6 la_data_in[17]
port 150 nsew default input
rlabel metal2 s 88191 0 88219 240 6 la_data_in[18]
port 151 nsew default input
rlabel metal2 s 89847 0 89875 240 6 la_data_in[19]
port 152 nsew default input
rlabel metal2 s 60177 0 60205 240 6 la_data_in[1]
port 153 nsew default input
rlabel metal2 s 91503 0 91531 240 6 la_data_in[20]
port 154 nsew default input
rlabel metal2 s 93159 0 93187 240 6 la_data_in[21]
port 155 nsew default input
rlabel metal2 s 94815 0 94843 240 6 la_data_in[22]
port 156 nsew default input
rlabel metal2 s 96471 0 96499 240 6 la_data_in[23]
port 157 nsew default input
rlabel metal2 s 98127 0 98155 240 6 la_data_in[24]
port 158 nsew default input
rlabel metal2 s 99737 0 99765 240 6 la_data_in[25]
port 159 nsew default input
rlabel metal2 s 101393 0 101421 240 6 la_data_in[26]
port 160 nsew default input
rlabel metal2 s 103049 0 103077 240 6 la_data_in[27]
port 161 nsew default input
rlabel metal2 s 104705 0 104733 240 6 la_data_in[28]
port 162 nsew default input
rlabel metal2 s 106361 0 106389 240 6 la_data_in[29]
port 163 nsew default input
rlabel metal2 s 61787 0 61815 240 6 la_data_in[2]
port 164 nsew default input
rlabel metal2 s 108017 0 108045 240 6 la_data_in[30]
port 165 nsew default input
rlabel metal2 s 109673 0 109701 240 6 la_data_in[31]
port 166 nsew default input
rlabel metal2 s 111283 0 111311 240 6 la_data_in[32]
port 167 nsew default input
rlabel metal2 s 112939 0 112967 240 6 la_data_in[33]
port 168 nsew default input
rlabel metal2 s 114595 0 114623 240 6 la_data_in[34]
port 169 nsew default input
rlabel metal2 s 116251 0 116279 240 6 la_data_in[35]
port 170 nsew default input
rlabel metal2 s 117907 0 117935 240 6 la_data_in[36]
port 171 nsew default input
rlabel metal2 s 119563 0 119591 240 6 la_data_in[37]
port 172 nsew default input
rlabel metal2 s 121219 0 121247 240 6 la_data_in[38]
port 173 nsew default input
rlabel metal2 s 122875 0 122903 240 6 la_data_in[39]
port 174 nsew default input
rlabel metal2 s 63443 0 63471 240 6 la_data_in[3]
port 175 nsew default input
rlabel metal2 s 124485 0 124513 240 6 la_data_in[40]
port 176 nsew default input
rlabel metal2 s 126141 0 126169 240 6 la_data_in[41]
port 177 nsew default input
rlabel metal2 s 127797 0 127825 240 6 la_data_in[42]
port 178 nsew default input
rlabel metal2 s 129453 0 129481 240 6 la_data_in[43]
port 179 nsew default input
rlabel metal2 s 131109 0 131137 240 6 la_data_in[44]
port 180 nsew default input
rlabel metal2 s 132765 0 132793 240 6 la_data_in[45]
port 181 nsew default input
rlabel metal2 s 134421 0 134449 240 6 la_data_in[46]
port 182 nsew default input
rlabel metal2 s 136031 0 136059 240 6 la_data_in[47]
port 183 nsew default input
rlabel metal2 s 137687 0 137715 240 6 la_data_in[48]
port 184 nsew default input
rlabel metal2 s 139343 0 139371 240 6 la_data_in[49]
port 185 nsew default input
rlabel metal2 s 65099 0 65127 240 6 la_data_in[4]
port 186 nsew default input
rlabel metal2 s 140999 0 141027 240 6 la_data_in[50]
port 187 nsew default input
rlabel metal2 s 142655 0 142683 240 6 la_data_in[51]
port 188 nsew default input
rlabel metal2 s 144311 0 144339 240 6 la_data_in[52]
port 189 nsew default input
rlabel metal2 s 145967 0 145995 240 6 la_data_in[53]
port 190 nsew default input
rlabel metal2 s 147577 0 147605 240 6 la_data_in[54]
port 191 nsew default input
rlabel metal2 s 149233 0 149261 240 6 la_data_in[55]
port 192 nsew default input
rlabel metal2 s 150889 0 150917 240 6 la_data_in[56]
port 193 nsew default input
rlabel metal2 s 152545 0 152573 240 6 la_data_in[57]
port 194 nsew default input
rlabel metal2 s 154201 0 154229 240 6 la_data_in[58]
port 195 nsew default input
rlabel metal2 s 155857 0 155885 240 6 la_data_in[59]
port 196 nsew default input
rlabel metal2 s 66755 0 66783 240 6 la_data_in[5]
port 197 nsew default input
rlabel metal2 s 157513 0 157541 240 6 la_data_in[60]
port 198 nsew default input
rlabel metal2 s 159169 0 159197 240 6 la_data_in[61]
port 199 nsew default input
rlabel metal2 s 160779 0 160807 240 6 la_data_in[62]
port 200 nsew default input
rlabel metal2 s 162435 0 162463 240 6 la_data_in[63]
port 201 nsew default input
rlabel metal2 s 164091 0 164119 240 6 la_data_in[64]
port 202 nsew default input
rlabel metal2 s 165747 0 165775 240 6 la_data_in[65]
port 203 nsew default input
rlabel metal2 s 167403 0 167431 240 6 la_data_in[66]
port 204 nsew default input
rlabel metal2 s 169059 0 169087 240 6 la_data_in[67]
port 205 nsew default input
rlabel metal2 s 170715 0 170743 240 6 la_data_in[68]
port 206 nsew default input
rlabel metal2 s 172325 0 172353 240 6 la_data_in[69]
port 207 nsew default input
rlabel metal2 s 68411 0 68439 240 6 la_data_in[6]
port 208 nsew default input
rlabel metal2 s 173981 0 174009 240 6 la_data_in[70]
port 209 nsew default input
rlabel metal2 s 175637 0 175665 240 6 la_data_in[71]
port 210 nsew default input
rlabel metal2 s 177293 0 177321 240 6 la_data_in[72]
port 211 nsew default input
rlabel metal2 s 178949 0 178977 240 6 la_data_in[73]
port 212 nsew default input
rlabel metal2 s 180605 0 180633 240 6 la_data_in[74]
port 213 nsew default input
rlabel metal2 s 182261 0 182289 240 6 la_data_in[75]
port 214 nsew default input
rlabel metal2 s 183917 0 183945 240 6 la_data_in[76]
port 215 nsew default input
rlabel metal2 s 185527 0 185555 240 6 la_data_in[77]
port 216 nsew default input
rlabel metal2 s 187183 0 187211 240 6 la_data_in[78]
port 217 nsew default input
rlabel metal2 s 188839 0 188867 240 6 la_data_in[79]
port 218 nsew default input
rlabel metal2 s 70067 0 70095 240 6 la_data_in[7]
port 219 nsew default input
rlabel metal2 s 190495 0 190523 240 6 la_data_in[80]
port 220 nsew default input
rlabel metal2 s 192151 0 192179 240 6 la_data_in[81]
port 221 nsew default input
rlabel metal2 s 193807 0 193835 240 6 la_data_in[82]
port 222 nsew default input
rlabel metal2 s 195463 0 195491 240 6 la_data_in[83]
port 223 nsew default input
rlabel metal2 s 197073 0 197101 240 6 la_data_in[84]
port 224 nsew default input
rlabel metal2 s 198729 0 198757 240 6 la_data_in[85]
port 225 nsew default input
rlabel metal2 s 200385 0 200413 240 6 la_data_in[86]
port 226 nsew default input
rlabel metal2 s 202041 0 202069 240 6 la_data_in[87]
port 227 nsew default input
rlabel metal2 s 203697 0 203725 240 6 la_data_in[88]
port 228 nsew default input
rlabel metal2 s 205353 0 205381 240 6 la_data_in[89]
port 229 nsew default input
rlabel metal2 s 71723 0 71751 240 6 la_data_in[8]
port 230 nsew default input
rlabel metal2 s 207009 0 207037 240 6 la_data_in[90]
port 231 nsew default input
rlabel metal2 s 208665 0 208693 240 6 la_data_in[91]
port 232 nsew default input
rlabel metal2 s 210275 0 210303 240 6 la_data_in[92]
port 233 nsew default input
rlabel metal2 s 211931 0 211959 240 6 la_data_in[93]
port 234 nsew default input
rlabel metal2 s 213587 0 213615 240 6 la_data_in[94]
port 235 nsew default input
rlabel metal2 s 215243 0 215271 240 6 la_data_in[95]
port 236 nsew default input
rlabel metal2 s 216899 0 216927 240 6 la_data_in[96]
port 237 nsew default input
rlabel metal2 s 218555 0 218583 240 6 la_data_in[97]
port 238 nsew default input
rlabel metal2 s 220211 0 220239 240 6 la_data_in[98]
port 239 nsew default input
rlabel metal2 s 221821 0 221849 240 6 la_data_in[99]
port 240 nsew default input
rlabel metal2 s 73379 0 73407 240 6 la_data_in[9]
port 241 nsew default input
rlabel metal2 s 59073 0 59101 240 6 la_data_out[0]
port 242 nsew default tristate
rlabel metal2 s 224029 0 224057 240 6 la_data_out[100]
port 243 nsew default tristate
rlabel metal2 s 225685 0 225713 240 6 la_data_out[101]
port 244 nsew default tristate
rlabel metal2 s 227341 0 227369 240 6 la_data_out[102]
port 245 nsew default tristate
rlabel metal2 s 228997 0 229025 240 6 la_data_out[103]
port 246 nsew default tristate
rlabel metal2 s 230653 0 230681 240 6 la_data_out[104]
port 247 nsew default tristate
rlabel metal2 s 232309 0 232337 240 6 la_data_out[105]
port 248 nsew default tristate
rlabel metal2 s 233919 0 233947 240 6 la_data_out[106]
port 249 nsew default tristate
rlabel metal2 s 235575 0 235603 240 6 la_data_out[107]
port 250 nsew default tristate
rlabel metal2 s 237231 0 237259 240 6 la_data_out[108]
port 251 nsew default tristate
rlabel metal2 s 238887 0 238915 240 6 la_data_out[109]
port 252 nsew default tristate
rlabel metal2 s 75541 0 75569 240 6 la_data_out[10]
port 253 nsew default tristate
rlabel metal2 s 240543 0 240571 240 6 la_data_out[110]
port 254 nsew default tristate
rlabel metal2 s 242199 0 242227 240 6 la_data_out[111]
port 255 nsew default tristate
rlabel metal2 s 243855 0 243883 240 6 la_data_out[112]
port 256 nsew default tristate
rlabel metal2 s 245511 0 245539 240 6 la_data_out[113]
port 257 nsew default tristate
rlabel metal2 s 247121 0 247149 240 6 la_data_out[114]
port 258 nsew default tristate
rlabel metal2 s 248777 0 248805 240 6 la_data_out[115]
port 259 nsew default tristate
rlabel metal2 s 250433 0 250461 240 6 la_data_out[116]
port 260 nsew default tristate
rlabel metal2 s 252089 0 252117 240 6 la_data_out[117]
port 261 nsew default tristate
rlabel metal2 s 253745 0 253773 240 6 la_data_out[118]
port 262 nsew default tristate
rlabel metal2 s 255401 0 255429 240 6 la_data_out[119]
port 263 nsew default tristate
rlabel metal2 s 77197 0 77225 240 6 la_data_out[11]
port 264 nsew default tristate
rlabel metal2 s 257057 0 257085 240 6 la_data_out[120]
port 265 nsew default tristate
rlabel metal2 s 258667 0 258695 240 6 la_data_out[121]
port 266 nsew default tristate
rlabel metal2 s 260323 0 260351 240 6 la_data_out[122]
port 267 nsew default tristate
rlabel metal2 s 261979 0 262007 240 6 la_data_out[123]
port 268 nsew default tristate
rlabel metal2 s 263635 0 263663 240 6 la_data_out[124]
port 269 nsew default tristate
rlabel metal2 s 265291 0 265319 240 6 la_data_out[125]
port 270 nsew default tristate
rlabel metal2 s 266947 0 266975 240 6 la_data_out[126]
port 271 nsew default tristate
rlabel metal2 s 268603 0 268631 240 6 la_data_out[127]
port 272 nsew default tristate
rlabel metal2 s 78853 0 78881 240 6 la_data_out[12]
port 273 nsew default tristate
rlabel metal2 s 80509 0 80537 240 6 la_data_out[13]
port 274 nsew default tristate
rlabel metal2 s 82165 0 82193 240 6 la_data_out[14]
port 275 nsew default tristate
rlabel metal2 s 83821 0 83849 240 6 la_data_out[15]
port 276 nsew default tristate
rlabel metal2 s 85477 0 85505 240 6 la_data_out[16]
port 277 nsew default tristate
rlabel metal2 s 87087 0 87115 240 6 la_data_out[17]
port 278 nsew default tristate
rlabel metal2 s 88743 0 88771 240 6 la_data_out[18]
port 279 nsew default tristate
rlabel metal2 s 90399 0 90427 240 6 la_data_out[19]
port 280 nsew default tristate
rlabel metal2 s 60729 0 60757 240 6 la_data_out[1]
port 281 nsew default tristate
rlabel metal2 s 92055 0 92083 240 6 la_data_out[20]
port 282 nsew default tristate
rlabel metal2 s 93711 0 93739 240 6 la_data_out[21]
port 283 nsew default tristate
rlabel metal2 s 95367 0 95395 240 6 la_data_out[22]
port 284 nsew default tristate
rlabel metal2 s 97023 0 97051 240 6 la_data_out[23]
port 285 nsew default tristate
rlabel metal2 s 98633 0 98661 240 6 la_data_out[24]
port 286 nsew default tristate
rlabel metal2 s 100289 0 100317 240 6 la_data_out[25]
port 287 nsew default tristate
rlabel metal2 s 101945 0 101973 240 6 la_data_out[26]
port 288 nsew default tristate
rlabel metal2 s 103601 0 103629 240 6 la_data_out[27]
port 289 nsew default tristate
rlabel metal2 s 105257 0 105285 240 6 la_data_out[28]
port 290 nsew default tristate
rlabel metal2 s 106913 0 106941 240 6 la_data_out[29]
port 291 nsew default tristate
rlabel metal2 s 62339 0 62367 240 6 la_data_out[2]
port 292 nsew default tristate
rlabel metal2 s 108569 0 108597 240 6 la_data_out[30]
port 293 nsew default tristate
rlabel metal2 s 110225 0 110253 240 6 la_data_out[31]
port 294 nsew default tristate
rlabel metal2 s 111835 0 111863 240 6 la_data_out[32]
port 295 nsew default tristate
rlabel metal2 s 113491 0 113519 240 6 la_data_out[33]
port 296 nsew default tristate
rlabel metal2 s 115147 0 115175 240 6 la_data_out[34]
port 297 nsew default tristate
rlabel metal2 s 116803 0 116831 240 6 la_data_out[35]
port 298 nsew default tristate
rlabel metal2 s 118459 0 118487 240 6 la_data_out[36]
port 299 nsew default tristate
rlabel metal2 s 120115 0 120143 240 6 la_data_out[37]
port 300 nsew default tristate
rlabel metal2 s 121771 0 121799 240 6 la_data_out[38]
port 301 nsew default tristate
rlabel metal2 s 123381 0 123409 240 6 la_data_out[39]
port 302 nsew default tristate
rlabel metal2 s 63995 0 64023 240 6 la_data_out[3]
port 303 nsew default tristate
rlabel metal2 s 125037 0 125065 240 6 la_data_out[40]
port 304 nsew default tristate
rlabel metal2 s 126693 0 126721 240 6 la_data_out[41]
port 305 nsew default tristate
rlabel metal2 s 128349 0 128377 240 6 la_data_out[42]
port 306 nsew default tristate
rlabel metal2 s 130005 0 130033 240 6 la_data_out[43]
port 307 nsew default tristate
rlabel metal2 s 131661 0 131689 240 6 la_data_out[44]
port 308 nsew default tristate
rlabel metal2 s 133317 0 133345 240 6 la_data_out[45]
port 309 nsew default tristate
rlabel metal2 s 134973 0 135001 240 6 la_data_out[46]
port 310 nsew default tristate
rlabel metal2 s 136583 0 136611 240 6 la_data_out[47]
port 311 nsew default tristate
rlabel metal2 s 138239 0 138267 240 6 la_data_out[48]
port 312 nsew default tristate
rlabel metal2 s 139895 0 139923 240 6 la_data_out[49]
port 313 nsew default tristate
rlabel metal2 s 65651 0 65679 240 6 la_data_out[4]
port 314 nsew default tristate
rlabel metal2 s 141551 0 141579 240 6 la_data_out[50]
port 315 nsew default tristate
rlabel metal2 s 143207 0 143235 240 6 la_data_out[51]
port 316 nsew default tristate
rlabel metal2 s 144863 0 144891 240 6 la_data_out[52]
port 317 nsew default tristate
rlabel metal2 s 146519 0 146547 240 6 la_data_out[53]
port 318 nsew default tristate
rlabel metal2 s 148129 0 148157 240 6 la_data_out[54]
port 319 nsew default tristate
rlabel metal2 s 149785 0 149813 240 6 la_data_out[55]
port 320 nsew default tristate
rlabel metal2 s 151441 0 151469 240 6 la_data_out[56]
port 321 nsew default tristate
rlabel metal2 s 153097 0 153125 240 6 la_data_out[57]
port 322 nsew default tristate
rlabel metal2 s 154753 0 154781 240 6 la_data_out[58]
port 323 nsew default tristate
rlabel metal2 s 156409 0 156437 240 6 la_data_out[59]
port 324 nsew default tristate
rlabel metal2 s 67307 0 67335 240 6 la_data_out[5]
port 325 nsew default tristate
rlabel metal2 s 158065 0 158093 240 6 la_data_out[60]
port 326 nsew default tristate
rlabel metal2 s 159721 0 159749 240 6 la_data_out[61]
port 327 nsew default tristate
rlabel metal2 s 161331 0 161359 240 6 la_data_out[62]
port 328 nsew default tristate
rlabel metal2 s 162987 0 163015 240 6 la_data_out[63]
port 329 nsew default tristate
rlabel metal2 s 164643 0 164671 240 6 la_data_out[64]
port 330 nsew default tristate
rlabel metal2 s 166299 0 166327 240 6 la_data_out[65]
port 331 nsew default tristate
rlabel metal2 s 167955 0 167983 240 6 la_data_out[66]
port 332 nsew default tristate
rlabel metal2 s 169611 0 169639 240 6 la_data_out[67]
port 333 nsew default tristate
rlabel metal2 s 171267 0 171295 240 6 la_data_out[68]
port 334 nsew default tristate
rlabel metal2 s 172877 0 172905 240 6 la_data_out[69]
port 335 nsew default tristate
rlabel metal2 s 68963 0 68991 240 6 la_data_out[6]
port 336 nsew default tristate
rlabel metal2 s 174533 0 174561 240 6 la_data_out[70]
port 337 nsew default tristate
rlabel metal2 s 176189 0 176217 240 6 la_data_out[71]
port 338 nsew default tristate
rlabel metal2 s 177845 0 177873 240 6 la_data_out[72]
port 339 nsew default tristate
rlabel metal2 s 179501 0 179529 240 6 la_data_out[73]
port 340 nsew default tristate
rlabel metal2 s 181157 0 181185 240 6 la_data_out[74]
port 341 nsew default tristate
rlabel metal2 s 182813 0 182841 240 6 la_data_out[75]
port 342 nsew default tristate
rlabel metal2 s 184423 0 184451 240 6 la_data_out[76]
port 343 nsew default tristate
rlabel metal2 s 186079 0 186107 240 6 la_data_out[77]
port 344 nsew default tristate
rlabel metal2 s 187735 0 187763 240 6 la_data_out[78]
port 345 nsew default tristate
rlabel metal2 s 189391 0 189419 240 6 la_data_out[79]
port 346 nsew default tristate
rlabel metal2 s 70619 0 70647 240 6 la_data_out[7]
port 347 nsew default tristate
rlabel metal2 s 191047 0 191075 240 6 la_data_out[80]
port 348 nsew default tristate
rlabel metal2 s 192703 0 192731 240 6 la_data_out[81]
port 349 nsew default tristate
rlabel metal2 s 194359 0 194387 240 6 la_data_out[82]
port 350 nsew default tristate
rlabel metal2 s 196015 0 196043 240 6 la_data_out[83]
port 351 nsew default tristate
rlabel metal2 s 197625 0 197653 240 6 la_data_out[84]
port 352 nsew default tristate
rlabel metal2 s 199281 0 199309 240 6 la_data_out[85]
port 353 nsew default tristate
rlabel metal2 s 200937 0 200965 240 6 la_data_out[86]
port 354 nsew default tristate
rlabel metal2 s 202593 0 202621 240 6 la_data_out[87]
port 355 nsew default tristate
rlabel metal2 s 204249 0 204277 240 6 la_data_out[88]
port 356 nsew default tristate
rlabel metal2 s 205905 0 205933 240 6 la_data_out[89]
port 357 nsew default tristate
rlabel metal2 s 72275 0 72303 240 6 la_data_out[8]
port 358 nsew default tristate
rlabel metal2 s 207561 0 207589 240 6 la_data_out[90]
port 359 nsew default tristate
rlabel metal2 s 209171 0 209199 240 6 la_data_out[91]
port 360 nsew default tristate
rlabel metal2 s 210827 0 210855 240 6 la_data_out[92]
port 361 nsew default tristate
rlabel metal2 s 212483 0 212511 240 6 la_data_out[93]
port 362 nsew default tristate
rlabel metal2 s 214139 0 214167 240 6 la_data_out[94]
port 363 nsew default tristate
rlabel metal2 s 215795 0 215823 240 6 la_data_out[95]
port 364 nsew default tristate
rlabel metal2 s 217451 0 217479 240 6 la_data_out[96]
port 365 nsew default tristate
rlabel metal2 s 219107 0 219135 240 6 la_data_out[97]
port 366 nsew default tristate
rlabel metal2 s 220763 0 220791 240 6 la_data_out[98]
port 367 nsew default tristate
rlabel metal2 s 222373 0 222401 240 6 la_data_out[99]
port 368 nsew default tristate
rlabel metal2 s 73885 0 73913 240 6 la_data_out[9]
port 369 nsew default tristate
rlabel metal2 s 59625 0 59653 240 6 la_oen[0]
port 370 nsew default input
rlabel metal2 s 224581 0 224609 240 6 la_oen[100]
port 371 nsew default input
rlabel metal2 s 226237 0 226265 240 6 la_oen[101]
port 372 nsew default input
rlabel metal2 s 227893 0 227921 240 6 la_oen[102]
port 373 nsew default input
rlabel metal2 s 229549 0 229577 240 6 la_oen[103]
port 374 nsew default input
rlabel metal2 s 231205 0 231233 240 6 la_oen[104]
port 375 nsew default input
rlabel metal2 s 232861 0 232889 240 6 la_oen[105]
port 376 nsew default input
rlabel metal2 s 234471 0 234499 240 6 la_oen[106]
port 377 nsew default input
rlabel metal2 s 236127 0 236155 240 6 la_oen[107]
port 378 nsew default input
rlabel metal2 s 237783 0 237811 240 6 la_oen[108]
port 379 nsew default input
rlabel metal2 s 239439 0 239467 240 6 la_oen[109]
port 380 nsew default input
rlabel metal2 s 76093 0 76121 240 6 la_oen[10]
port 381 nsew default input
rlabel metal2 s 241095 0 241123 240 6 la_oen[110]
port 382 nsew default input
rlabel metal2 s 242751 0 242779 240 6 la_oen[111]
port 383 nsew default input
rlabel metal2 s 244407 0 244435 240 6 la_oen[112]
port 384 nsew default input
rlabel metal2 s 246017 0 246045 240 6 la_oen[113]
port 385 nsew default input
rlabel metal2 s 247673 0 247701 240 6 la_oen[114]
port 386 nsew default input
rlabel metal2 s 249329 0 249357 240 6 la_oen[115]
port 387 nsew default input
rlabel metal2 s 250985 0 251013 240 6 la_oen[116]
port 388 nsew default input
rlabel metal2 s 252641 0 252669 240 6 la_oen[117]
port 389 nsew default input
rlabel metal2 s 254297 0 254325 240 6 la_oen[118]
port 390 nsew default input
rlabel metal2 s 255953 0 255981 240 6 la_oen[119]
port 391 nsew default input
rlabel metal2 s 77749 0 77777 240 6 la_oen[11]
port 392 nsew default input
rlabel metal2 s 257609 0 257637 240 6 la_oen[120]
port 393 nsew default input
rlabel metal2 s 259219 0 259247 240 6 la_oen[121]
port 394 nsew default input
rlabel metal2 s 260875 0 260903 240 6 la_oen[122]
port 395 nsew default input
rlabel metal2 s 262531 0 262559 240 6 la_oen[123]
port 396 nsew default input
rlabel metal2 s 264187 0 264215 240 6 la_oen[124]
port 397 nsew default input
rlabel metal2 s 265843 0 265871 240 6 la_oen[125]
port 398 nsew default input
rlabel metal2 s 267499 0 267527 240 6 la_oen[126]
port 399 nsew default input
rlabel metal2 s 269155 0 269183 240 6 la_oen[127]
port 400 nsew default input
rlabel metal2 s 79405 0 79433 240 6 la_oen[12]
port 401 nsew default input
rlabel metal2 s 81061 0 81089 240 6 la_oen[13]
port 402 nsew default input
rlabel metal2 s 82717 0 82745 240 6 la_oen[14]
port 403 nsew default input
rlabel metal2 s 84373 0 84401 240 6 la_oen[15]
port 404 nsew default input
rlabel metal2 s 86029 0 86057 240 6 la_oen[16]
port 405 nsew default input
rlabel metal2 s 87639 0 87667 240 6 la_oen[17]
port 406 nsew default input
rlabel metal2 s 89295 0 89323 240 6 la_oen[18]
port 407 nsew default input
rlabel metal2 s 90951 0 90979 240 6 la_oen[19]
port 408 nsew default input
rlabel metal2 s 61281 0 61309 240 6 la_oen[1]
port 409 nsew default input
rlabel metal2 s 92607 0 92635 240 6 la_oen[20]
port 410 nsew default input
rlabel metal2 s 94263 0 94291 240 6 la_oen[21]
port 411 nsew default input
rlabel metal2 s 95919 0 95947 240 6 la_oen[22]
port 412 nsew default input
rlabel metal2 s 97575 0 97603 240 6 la_oen[23]
port 413 nsew default input
rlabel metal2 s 99185 0 99213 240 6 la_oen[24]
port 414 nsew default input
rlabel metal2 s 100841 0 100869 240 6 la_oen[25]
port 415 nsew default input
rlabel metal2 s 102497 0 102525 240 6 la_oen[26]
port 416 nsew default input
rlabel metal2 s 104153 0 104181 240 6 la_oen[27]
port 417 nsew default input
rlabel metal2 s 105809 0 105837 240 6 la_oen[28]
port 418 nsew default input
rlabel metal2 s 107465 0 107493 240 6 la_oen[29]
port 419 nsew default input
rlabel metal2 s 62891 0 62919 240 6 la_oen[2]
port 420 nsew default input
rlabel metal2 s 109121 0 109149 240 6 la_oen[30]
port 421 nsew default input
rlabel metal2 s 110731 0 110759 240 6 la_oen[31]
port 422 nsew default input
rlabel metal2 s 112387 0 112415 240 6 la_oen[32]
port 423 nsew default input
rlabel metal2 s 114043 0 114071 240 6 la_oen[33]
port 424 nsew default input
rlabel metal2 s 115699 0 115727 240 6 la_oen[34]
port 425 nsew default input
rlabel metal2 s 117355 0 117383 240 6 la_oen[35]
port 426 nsew default input
rlabel metal2 s 119011 0 119039 240 6 la_oen[36]
port 427 nsew default input
rlabel metal2 s 120667 0 120695 240 6 la_oen[37]
port 428 nsew default input
rlabel metal2 s 122323 0 122351 240 6 la_oen[38]
port 429 nsew default input
rlabel metal2 s 123933 0 123961 240 6 la_oen[39]
port 430 nsew default input
rlabel metal2 s 64547 0 64575 240 6 la_oen[3]
port 431 nsew default input
rlabel metal2 s 125589 0 125617 240 6 la_oen[40]
port 432 nsew default input
rlabel metal2 s 127245 0 127273 240 6 la_oen[41]
port 433 nsew default input
rlabel metal2 s 128901 0 128929 240 6 la_oen[42]
port 434 nsew default input
rlabel metal2 s 130557 0 130585 240 6 la_oen[43]
port 435 nsew default input
rlabel metal2 s 132213 0 132241 240 6 la_oen[44]
port 436 nsew default input
rlabel metal2 s 133869 0 133897 240 6 la_oen[45]
port 437 nsew default input
rlabel metal2 s 135479 0 135507 240 6 la_oen[46]
port 438 nsew default input
rlabel metal2 s 137135 0 137163 240 6 la_oen[47]
port 439 nsew default input
rlabel metal2 s 138791 0 138819 240 6 la_oen[48]
port 440 nsew default input
rlabel metal2 s 140447 0 140475 240 6 la_oen[49]
port 441 nsew default input
rlabel metal2 s 66203 0 66231 240 6 la_oen[4]
port 442 nsew default input
rlabel metal2 s 142103 0 142131 240 6 la_oen[50]
port 443 nsew default input
rlabel metal2 s 143759 0 143787 240 6 la_oen[51]
port 444 nsew default input
rlabel metal2 s 145415 0 145443 240 6 la_oen[52]
port 445 nsew default input
rlabel metal2 s 147071 0 147099 240 6 la_oen[53]
port 446 nsew default input
rlabel metal2 s 148681 0 148709 240 6 la_oen[54]
port 447 nsew default input
rlabel metal2 s 150337 0 150365 240 6 la_oen[55]
port 448 nsew default input
rlabel metal2 s 151993 0 152021 240 6 la_oen[56]
port 449 nsew default input
rlabel metal2 s 153649 0 153677 240 6 la_oen[57]
port 450 nsew default input
rlabel metal2 s 155305 0 155333 240 6 la_oen[58]
port 451 nsew default input
rlabel metal2 s 156961 0 156989 240 6 la_oen[59]
port 452 nsew default input
rlabel metal2 s 67859 0 67887 240 6 la_oen[5]
port 453 nsew default input
rlabel metal2 s 158617 0 158645 240 6 la_oen[60]
port 454 nsew default input
rlabel metal2 s 160227 0 160255 240 6 la_oen[61]
port 455 nsew default input
rlabel metal2 s 161883 0 161911 240 6 la_oen[62]
port 456 nsew default input
rlabel metal2 s 163539 0 163567 240 6 la_oen[63]
port 457 nsew default input
rlabel metal2 s 165195 0 165223 240 6 la_oen[64]
port 458 nsew default input
rlabel metal2 s 166851 0 166879 240 6 la_oen[65]
port 459 nsew default input
rlabel metal2 s 168507 0 168535 240 6 la_oen[66]
port 460 nsew default input
rlabel metal2 s 170163 0 170191 240 6 la_oen[67]
port 461 nsew default input
rlabel metal2 s 171819 0 171847 240 6 la_oen[68]
port 462 nsew default input
rlabel metal2 s 173429 0 173457 240 6 la_oen[69]
port 463 nsew default input
rlabel metal2 s 69515 0 69543 240 6 la_oen[6]
port 464 nsew default input
rlabel metal2 s 175085 0 175113 240 6 la_oen[70]
port 465 nsew default input
rlabel metal2 s 176741 0 176769 240 6 la_oen[71]
port 466 nsew default input
rlabel metal2 s 178397 0 178425 240 6 la_oen[72]
port 467 nsew default input
rlabel metal2 s 180053 0 180081 240 6 la_oen[73]
port 468 nsew default input
rlabel metal2 s 181709 0 181737 240 6 la_oen[74]
port 469 nsew default input
rlabel metal2 s 183365 0 183393 240 6 la_oen[75]
port 470 nsew default input
rlabel metal2 s 184975 0 185003 240 6 la_oen[76]
port 471 nsew default input
rlabel metal2 s 186631 0 186659 240 6 la_oen[77]
port 472 nsew default input
rlabel metal2 s 188287 0 188315 240 6 la_oen[78]
port 473 nsew default input
rlabel metal2 s 189943 0 189971 240 6 la_oen[79]
port 474 nsew default input
rlabel metal2 s 71171 0 71199 240 6 la_oen[7]
port 475 nsew default input
rlabel metal2 s 191599 0 191627 240 6 la_oen[80]
port 476 nsew default input
rlabel metal2 s 193255 0 193283 240 6 la_oen[81]
port 477 nsew default input
rlabel metal2 s 194911 0 194939 240 6 la_oen[82]
port 478 nsew default input
rlabel metal2 s 196567 0 196595 240 6 la_oen[83]
port 479 nsew default input
rlabel metal2 s 198177 0 198205 240 6 la_oen[84]
port 480 nsew default input
rlabel metal2 s 199833 0 199861 240 6 la_oen[85]
port 481 nsew default input
rlabel metal2 s 201489 0 201517 240 6 la_oen[86]
port 482 nsew default input
rlabel metal2 s 203145 0 203173 240 6 la_oen[87]
port 483 nsew default input
rlabel metal2 s 204801 0 204829 240 6 la_oen[88]
port 484 nsew default input
rlabel metal2 s 206457 0 206485 240 6 la_oen[89]
port 485 nsew default input
rlabel metal2 s 72827 0 72855 240 6 la_oen[8]
port 486 nsew default input
rlabel metal2 s 208113 0 208141 240 6 la_oen[90]
port 487 nsew default input
rlabel metal2 s 209723 0 209751 240 6 la_oen[91]
port 488 nsew default input
rlabel metal2 s 211379 0 211407 240 6 la_oen[92]
port 489 nsew default input
rlabel metal2 s 213035 0 213063 240 6 la_oen[93]
port 490 nsew default input
rlabel metal2 s 214691 0 214719 240 6 la_oen[94]
port 491 nsew default input
rlabel metal2 s 216347 0 216375 240 6 la_oen[95]
port 492 nsew default input
rlabel metal2 s 218003 0 218031 240 6 la_oen[96]
port 493 nsew default input
rlabel metal2 s 219659 0 219687 240 6 la_oen[97]
port 494 nsew default input
rlabel metal2 s 221269 0 221297 240 6 la_oen[98]
port 495 nsew default input
rlabel metal2 s 222925 0 222953 240 6 la_oen[99]
port 496 nsew default input
rlabel metal2 s 74437 0 74465 240 6 la_oen[9]
port 497 nsew default input
rlabel metal2 s 269707 0 269735 240 6 user_clock2
port 498 nsew default input
rlabel metal3 s 269760 250312 270000 250372 6 vccd1
port 499 nsew default bidirectional
rlabel metal3 s 0 249428 240 249488 6 vccd2
port 500 nsew default bidirectional
rlabel metal3 s 269760 126552 270000 126612 6 vdda1
port 501 nsew default bidirectional
rlabel metal3 s 0 114448 240 114508 6 vdda2
port 502 nsew default bidirectional
rlabel metal2 s 236219 269760 236247 270000 6 vssa1
port 503 nsew default bidirectional
rlabel metal3 s 0 243580 240 243640 6 vssa2
port 504 nsew default bidirectional
rlabel metal3 s 269760 120908 270000 120968 6 vssd1
port 505 nsew default bidirectional
rlabel metal3 s 0 108532 240 108592 6 vssd2
port 506 nsew default bidirectional
rlabel metal2 s 239 0 267 240 6 wb_clk_i
port 507 nsew default input
rlabel metal2 s 745 0 773 240 6 wb_rst_i
port 508 nsew default input
rlabel metal2 s 1297 0 1325 240 6 wbs_ack_o
port 509 nsew default tristate
rlabel metal2 s 3505 0 3533 240 6 wbs_adr_i[0]
port 510 nsew default input
rlabel metal2 s 22227 0 22255 240 6 wbs_adr_i[10]
port 511 nsew default input
rlabel metal2 s 23883 0 23911 240 6 wbs_adr_i[11]
port 512 nsew default input
rlabel metal2 s 25493 0 25521 240 6 wbs_adr_i[12]
port 513 nsew default input
rlabel metal2 s 27149 0 27177 240 6 wbs_adr_i[13]
port 514 nsew default input
rlabel metal2 s 28805 0 28833 240 6 wbs_adr_i[14]
port 515 nsew default input
rlabel metal2 s 30461 0 30489 240 6 wbs_adr_i[15]
port 516 nsew default input
rlabel metal2 s 32117 0 32145 240 6 wbs_adr_i[16]
port 517 nsew default input
rlabel metal2 s 33773 0 33801 240 6 wbs_adr_i[17]
port 518 nsew default input
rlabel metal2 s 35429 0 35457 240 6 wbs_adr_i[18]
port 519 nsew default input
rlabel metal2 s 37039 0 37067 240 6 wbs_adr_i[19]
port 520 nsew default input
rlabel metal2 s 5713 0 5741 240 6 wbs_adr_i[1]
port 521 nsew default input
rlabel metal2 s 38695 0 38723 240 6 wbs_adr_i[20]
port 522 nsew default input
rlabel metal2 s 40351 0 40379 240 6 wbs_adr_i[21]
port 523 nsew default input
rlabel metal2 s 42007 0 42035 240 6 wbs_adr_i[22]
port 524 nsew default input
rlabel metal2 s 43663 0 43691 240 6 wbs_adr_i[23]
port 525 nsew default input
rlabel metal2 s 45319 0 45347 240 6 wbs_adr_i[24]
port 526 nsew default input
rlabel metal2 s 46975 0 47003 240 6 wbs_adr_i[25]
port 527 nsew default input
rlabel metal2 s 48631 0 48659 240 6 wbs_adr_i[26]
port 528 nsew default input
rlabel metal2 s 50241 0 50269 240 6 wbs_adr_i[27]
port 529 nsew default input
rlabel metal2 s 51897 0 51925 240 6 wbs_adr_i[28]
port 530 nsew default input
rlabel metal2 s 53553 0 53581 240 6 wbs_adr_i[29]
port 531 nsew default input
rlabel metal2 s 7921 0 7949 240 6 wbs_adr_i[2]
port 532 nsew default input
rlabel metal2 s 55209 0 55237 240 6 wbs_adr_i[30]
port 533 nsew default input
rlabel metal2 s 56865 0 56893 240 6 wbs_adr_i[31]
port 534 nsew default input
rlabel metal2 s 10129 0 10157 240 6 wbs_adr_i[3]
port 535 nsew default input
rlabel metal2 s 12337 0 12365 240 6 wbs_adr_i[4]
port 536 nsew default input
rlabel metal2 s 13947 0 13975 240 6 wbs_adr_i[5]
port 537 nsew default input
rlabel metal2 s 15603 0 15631 240 6 wbs_adr_i[6]
port 538 nsew default input
rlabel metal2 s 17259 0 17287 240 6 wbs_adr_i[7]
port 539 nsew default input
rlabel metal2 s 18915 0 18943 240 6 wbs_adr_i[8]
port 540 nsew default input
rlabel metal2 s 20571 0 20599 240 6 wbs_adr_i[9]
port 541 nsew default input
rlabel metal2 s 1849 0 1877 240 6 wbs_cyc_i
port 542 nsew default input
rlabel metal2 s 4057 0 4085 240 6 wbs_dat_i[0]
port 543 nsew default input
rlabel metal2 s 22779 0 22807 240 6 wbs_dat_i[10]
port 544 nsew default input
rlabel metal2 s 24435 0 24463 240 6 wbs_dat_i[11]
port 545 nsew default input
rlabel metal2 s 26045 0 26073 240 6 wbs_dat_i[12]
port 546 nsew default input
rlabel metal2 s 27701 0 27729 240 6 wbs_dat_i[13]
port 547 nsew default input
rlabel metal2 s 29357 0 29385 240 6 wbs_dat_i[14]
port 548 nsew default input
rlabel metal2 s 31013 0 31041 240 6 wbs_dat_i[15]
port 549 nsew default input
rlabel metal2 s 32669 0 32697 240 6 wbs_dat_i[16]
port 550 nsew default input
rlabel metal2 s 34325 0 34353 240 6 wbs_dat_i[17]
port 551 nsew default input
rlabel metal2 s 35981 0 36009 240 6 wbs_dat_i[18]
port 552 nsew default input
rlabel metal2 s 37591 0 37619 240 6 wbs_dat_i[19]
port 553 nsew default input
rlabel metal2 s 6265 0 6293 240 6 wbs_dat_i[1]
port 554 nsew default input
rlabel metal2 s 39247 0 39275 240 6 wbs_dat_i[20]
port 555 nsew default input
rlabel metal2 s 40903 0 40931 240 6 wbs_dat_i[21]
port 556 nsew default input
rlabel metal2 s 42559 0 42587 240 6 wbs_dat_i[22]
port 557 nsew default input
rlabel metal2 s 44215 0 44243 240 6 wbs_dat_i[23]
port 558 nsew default input
rlabel metal2 s 45871 0 45899 240 6 wbs_dat_i[24]
port 559 nsew default input
rlabel metal2 s 47527 0 47555 240 6 wbs_dat_i[25]
port 560 nsew default input
rlabel metal2 s 49183 0 49211 240 6 wbs_dat_i[26]
port 561 nsew default input
rlabel metal2 s 50793 0 50821 240 6 wbs_dat_i[27]
port 562 nsew default input
rlabel metal2 s 52449 0 52477 240 6 wbs_dat_i[28]
port 563 nsew default input
rlabel metal2 s 54105 0 54133 240 6 wbs_dat_i[29]
port 564 nsew default input
rlabel metal2 s 8473 0 8501 240 6 wbs_dat_i[2]
port 565 nsew default input
rlabel metal2 s 55761 0 55789 240 6 wbs_dat_i[30]
port 566 nsew default input
rlabel metal2 s 57417 0 57445 240 6 wbs_dat_i[31]
port 567 nsew default input
rlabel metal2 s 10681 0 10709 240 6 wbs_dat_i[3]
port 568 nsew default input
rlabel metal2 s 12843 0 12871 240 6 wbs_dat_i[4]
port 569 nsew default input
rlabel metal2 s 14499 0 14527 240 6 wbs_dat_i[5]
port 570 nsew default input
rlabel metal2 s 16155 0 16183 240 6 wbs_dat_i[6]
port 571 nsew default input
rlabel metal2 s 17811 0 17839 240 6 wbs_dat_i[7]
port 572 nsew default input
rlabel metal2 s 19467 0 19495 240 6 wbs_dat_i[8]
port 573 nsew default input
rlabel metal2 s 21123 0 21151 240 6 wbs_dat_i[9]
port 574 nsew default input
rlabel metal2 s 4609 0 4637 240 6 wbs_dat_o[0]
port 575 nsew default tristate
rlabel metal2 s 23331 0 23359 240 6 wbs_dat_o[10]
port 576 nsew default tristate
rlabel metal2 s 24941 0 24969 240 6 wbs_dat_o[11]
port 577 nsew default tristate
rlabel metal2 s 26597 0 26625 240 6 wbs_dat_o[12]
port 578 nsew default tristate
rlabel metal2 s 28253 0 28281 240 6 wbs_dat_o[13]
port 579 nsew default tristate
rlabel metal2 s 29909 0 29937 240 6 wbs_dat_o[14]
port 580 nsew default tristate
rlabel metal2 s 31565 0 31593 240 6 wbs_dat_o[15]
port 581 nsew default tristate
rlabel metal2 s 33221 0 33249 240 6 wbs_dat_o[16]
port 582 nsew default tristate
rlabel metal2 s 34877 0 34905 240 6 wbs_dat_o[17]
port 583 nsew default tristate
rlabel metal2 s 36533 0 36561 240 6 wbs_dat_o[18]
port 584 nsew default tristate
rlabel metal2 s 38143 0 38171 240 6 wbs_dat_o[19]
port 585 nsew default tristate
rlabel metal2 s 6817 0 6845 240 6 wbs_dat_o[1]
port 586 nsew default tristate
rlabel metal2 s 39799 0 39827 240 6 wbs_dat_o[20]
port 587 nsew default tristate
rlabel metal2 s 41455 0 41483 240 6 wbs_dat_o[21]
port 588 nsew default tristate
rlabel metal2 s 43111 0 43139 240 6 wbs_dat_o[22]
port 589 nsew default tristate
rlabel metal2 s 44767 0 44795 240 6 wbs_dat_o[23]
port 590 nsew default tristate
rlabel metal2 s 46423 0 46451 240 6 wbs_dat_o[24]
port 591 nsew default tristate
rlabel metal2 s 48079 0 48107 240 6 wbs_dat_o[25]
port 592 nsew default tristate
rlabel metal2 s 49689 0 49717 240 6 wbs_dat_o[26]
port 593 nsew default tristate
rlabel metal2 s 51345 0 51373 240 6 wbs_dat_o[27]
port 594 nsew default tristate
rlabel metal2 s 53001 0 53029 240 6 wbs_dat_o[28]
port 595 nsew default tristate
rlabel metal2 s 54657 0 54685 240 6 wbs_dat_o[29]
port 596 nsew default tristate
rlabel metal2 s 9025 0 9053 240 6 wbs_dat_o[2]
port 597 nsew default tristate
rlabel metal2 s 56313 0 56341 240 6 wbs_dat_o[30]
port 598 nsew default tristate
rlabel metal2 s 57969 0 57997 240 6 wbs_dat_o[31]
port 599 nsew default tristate
rlabel metal2 s 11233 0 11261 240 6 wbs_dat_o[3]
port 600 nsew default tristate
rlabel metal2 s 13395 0 13423 240 6 wbs_dat_o[4]
port 601 nsew default tristate
rlabel metal2 s 15051 0 15079 240 6 wbs_dat_o[5]
port 602 nsew default tristate
rlabel metal2 s 16707 0 16735 240 6 wbs_dat_o[6]
port 603 nsew default tristate
rlabel metal2 s 18363 0 18391 240 6 wbs_dat_o[7]
port 604 nsew default tristate
rlabel metal2 s 20019 0 20047 240 6 wbs_dat_o[8]
port 605 nsew default tristate
rlabel metal2 s 21675 0 21703 240 6 wbs_dat_o[9]
port 606 nsew default tristate
rlabel metal2 s 5161 0 5189 240 6 wbs_sel_i[0]
port 607 nsew default input
rlabel metal2 s 7369 0 7397 240 6 wbs_sel_i[1]
port 608 nsew default input
rlabel metal2 s 9577 0 9605 240 6 wbs_sel_i[2]
port 609 nsew default input
rlabel metal2 s 11785 0 11813 240 6 wbs_sel_i[3]
port 610 nsew default input
rlabel metal2 s 2401 0 2429 240 6 wbs_stb_i
port 611 nsew default input
rlabel metal2 s 2953 0 2981 240 6 wbs_we_i
port 612 nsew default input
<< end >>
